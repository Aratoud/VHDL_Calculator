library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity shift_rpn_registers_down is
  Port 
  (
  );
end shift_rpn_registers_down;

architecture Behavioral of shift_rpn_registers_down is

begin


end Behavioral;

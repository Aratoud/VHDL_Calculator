library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity stringROM is
  Port 
  (
    reg0_int : in integer;
    reg1_int : in integer;
    reg2_int : in integer;
    reg3_int : in integer;
    
    reg0_string : out string(1 to 4);
    reg1_string : out string(1 to 4); 
    reg2_string : out string(1 to 4);
    reg3_string : out string(1 to 4) 
  );
end stringROM;

architecture Behavioral of stringROM is

begin

    reg0_LUT : process(reg3_int, reg2_int, reg1_int, reg0_int) 
    begin 
        case (reg3_int) is
            when 999 => reg3_string <= " 999";
            when 998 => reg3_string <= " 998";
            when 997 => reg3_string <= " 997";
            when 996 => reg3_string <= " 996";
            when 995 => reg3_string <= " 995";
            when 994 => reg3_string <= " 994";
            when 993 => reg3_string <= " 993";
            when 992 => reg3_string <= " 992";
            when 991 => reg3_string <= " 991";
            when 990 => reg3_string <= " 990";
            when 989 => reg3_string <= " 989";
            when 988 => reg3_string <= " 988";
            when 987 => reg3_string <= " 987";
            when 986 => reg3_string <= " 986";
            when 985 => reg3_string <= " 985";
            when 984 => reg3_string <= " 984";
            when 983 => reg3_string <= " 983";
            when 982 => reg3_string <= " 982";
            when 981 => reg3_string <= " 981";
            when 980 => reg3_string <= " 980";
            when 979 => reg3_string <= " 979";
            when 978 => reg3_string <= " 978";
            when 977 => reg3_string <= " 977";
            when 976 => reg3_string <= " 976";
            when 975 => reg3_string <= " 975";
            when 974 => reg3_string <= " 974";
            when 973 => reg3_string <= " 973";
            when 972 => reg3_string <= " 972";
            when 971 => reg3_string <= " 971";
            when 970 => reg3_string <= " 970";
            when 969 => reg3_string <= " 969";
            when 968 => reg3_string <= " 968";
            when 967 => reg3_string <= " 967";
            when 966 => reg3_string <= " 966";
            when 965 => reg3_string <= " 965";
            when 964 => reg3_string <= " 964";
            when 963 => reg3_string <= " 963";
            when 962 => reg3_string <= " 962";
            when 961 => reg3_string <= " 961";
            when 960 => reg3_string <= " 960";
            when 959 => reg3_string <= " 959";
            when 958 => reg3_string <= " 958";
            when 957 => reg3_string <= " 957";
            when 956 => reg3_string <= " 956";
            when 955 => reg3_string <= " 955";
            when 954 => reg3_string <= " 954";
            when 953 => reg3_string <= " 953";
            when 952 => reg3_string <= " 952";
            when 951 => reg3_string <= " 951";
            when 950 => reg3_string <= " 950";
            when 949 => reg3_string <= " 949";
            when 948 => reg3_string <= " 948";
            when 947 => reg3_string <= " 947";
            when 946 => reg3_string <= " 946";
            when 945 => reg3_string <= " 945";
            when 944 => reg3_string <= " 944";
            when 943 => reg3_string <= " 943";
            when 942 => reg3_string <= " 942";
            when 941 => reg3_string <= " 941";
            when 940 => reg3_string <= " 940";
            when 939 => reg3_string <= " 939";
            when 938 => reg3_string <= " 938";
            when 937 => reg3_string <= " 937";
            when 936 => reg3_string <= " 936";
            when 935 => reg3_string <= " 935";
            when 934 => reg3_string <= " 934";
            when 933 => reg3_string <= " 933";
            when 932 => reg3_string <= " 932";
            when 931 => reg3_string <= " 931";
            when 930 => reg3_string <= " 930";
            when 929 => reg3_string <= " 929";
            when 928 => reg3_string <= " 928";
            when 927 => reg3_string <= " 927";
            when 926 => reg3_string <= " 926";
            when 925 => reg3_string <= " 925";
            when 924 => reg3_string <= " 924";
            when 923 => reg3_string <= " 923";
            when 922 => reg3_string <= " 922";
            when 921 => reg3_string <= " 921";
            when 920 => reg3_string <= " 920";
            when 919 => reg3_string <= " 919";
            when 918 => reg3_string <= " 918";
            when 917 => reg3_string <= " 917";
            when 916 => reg3_string <= " 916";
            when 915 => reg3_string <= " 915";
            when 914 => reg3_string <= " 914";
            when 913 => reg3_string <= " 913";
            when 912 => reg3_string <= " 912";
            when 911 => reg3_string <= " 911";
            when 910 => reg3_string <= " 910";
            when 909 => reg3_string <= " 909";
            when 908 => reg3_string <= " 908";
            when 907 => reg3_string <= " 907";
            when 906 => reg3_string <= " 906";
            when 905 => reg3_string <= " 905";
            when 904 => reg3_string <= " 904";
            when 903 => reg3_string <= " 903";
            when 902 => reg3_string <= " 902";
            when 901 => reg3_string <= " 901";
            when 900 => reg3_string <= " 900";
            when 899 => reg3_string <= " 899";
            when 898 => reg3_string <= " 898";
            when 897 => reg3_string <= " 897";
            when 896 => reg3_string <= " 896";
            when 895 => reg3_string <= " 895";
            when 894 => reg3_string <= " 894";
            when 893 => reg3_string <= " 893";
            when 892 => reg3_string <= " 892";
            when 891 => reg3_string <= " 891";
            when 890 => reg3_string <= " 890";
            when 889 => reg3_string <= " 889";
            when 888 => reg3_string <= " 888";
            when 887 => reg3_string <= " 887";
            when 886 => reg3_string <= " 886";
            when 885 => reg3_string <= " 885";
            when 884 => reg3_string <= " 884";
            when 883 => reg3_string <= " 883";
            when 882 => reg3_string <= " 882";
            when 881 => reg3_string <= " 881";
            when 880 => reg3_string <= " 880";
            when 879 => reg3_string <= " 879";
            when 878 => reg3_string <= " 878";
            when 877 => reg3_string <= " 877";
            when 876 => reg3_string <= " 876";
            when 875 => reg3_string <= " 875";
            when 874 => reg3_string <= " 874";
            when 873 => reg3_string <= " 873";
            when 872 => reg3_string <= " 872";
            when 871 => reg3_string <= " 871";
            when 870 => reg3_string <= " 870";
            when 869 => reg3_string <= " 869";
            when 868 => reg3_string <= " 868";
            when 867 => reg3_string <= " 867";
            when 866 => reg3_string <= " 866";
            when 865 => reg3_string <= " 865";
            when 864 => reg3_string <= " 864";
            when 863 => reg3_string <= " 863";
            when 862 => reg3_string <= " 862";
            when 861 => reg3_string <= " 861";
            when 860 => reg3_string <= " 860";
            when 859 => reg3_string <= " 859";
            when 858 => reg3_string <= " 858";
            when 857 => reg3_string <= " 857";
            when 856 => reg3_string <= " 856";
            when 855 => reg3_string <= " 855";
            when 854 => reg3_string <= " 854";
            when 853 => reg3_string <= " 853";
            when 852 => reg3_string <= " 852";
            when 851 => reg3_string <= " 851";
            when 850 => reg3_string <= " 850";
            when 849 => reg3_string <= " 849";
            when 848 => reg3_string <= " 848";
            when 847 => reg3_string <= " 847";
            when 846 => reg3_string <= " 846";
            when 845 => reg3_string <= " 845";
            when 844 => reg3_string <= " 844";
            when 843 => reg3_string <= " 843";
            when 842 => reg3_string <= " 842";
            when 841 => reg3_string <= " 841";
            when 840 => reg3_string <= " 840";
            when 839 => reg3_string <= " 839";
            when 838 => reg3_string <= " 838";
            when 837 => reg3_string <= " 837";
            when 836 => reg3_string <= " 836";
            when 835 => reg3_string <= " 835";
            when 834 => reg3_string <= " 834";
            when 833 => reg3_string <= " 833";
            when 832 => reg3_string <= " 832";
            when 831 => reg3_string <= " 831";
            when 830 => reg3_string <= " 830";
            when 829 => reg3_string <= " 829";
            when 828 => reg3_string <= " 828";
            when 827 => reg3_string <= " 827";
            when 826 => reg3_string <= " 826";
            when 825 => reg3_string <= " 825";
            when 824 => reg3_string <= " 824";
            when 823 => reg3_string <= " 823";
            when 822 => reg3_string <= " 822";
            when 821 => reg3_string <= " 821";
            when 820 => reg3_string <= " 820";
            when 819 => reg3_string <= " 819";
            when 818 => reg3_string <= " 818";
            when 817 => reg3_string <= " 817";
            when 816 => reg3_string <= " 816";
            when 815 => reg3_string <= " 815";
            when 814 => reg3_string <= " 814";
            when 813 => reg3_string <= " 813";
            when 812 => reg3_string <= " 812";
            when 811 => reg3_string <= " 811";
            when 810 => reg3_string <= " 810";
            when 809 => reg3_string <= " 809";
            when 808 => reg3_string <= " 808";
            when 807 => reg3_string <= " 807";
            when 806 => reg3_string <= " 806";
            when 805 => reg3_string <= " 805";
            when 804 => reg3_string <= " 804";
            when 803 => reg3_string <= " 803";
            when 802 => reg3_string <= " 802";
            when 801 => reg3_string <= " 801";
            when 800 => reg3_string <= " 800";
            when 799 => reg3_string <= " 799";
            when 798 => reg3_string <= " 798";
            when 797 => reg3_string <= " 797";
            when 796 => reg3_string <= " 796";
            when 795 => reg3_string <= " 795";
            when 794 => reg3_string <= " 794";
            when 793 => reg3_string <= " 793";
            when 792 => reg3_string <= " 792";
            when 791 => reg3_string <= " 791";
            when 790 => reg3_string <= " 790";
            when 789 => reg3_string <= " 789";
            when 788 => reg3_string <= " 788";
            when 787 => reg3_string <= " 787";
            when 786 => reg3_string <= " 786";
            when 785 => reg3_string <= " 785";
            when 784 => reg3_string <= " 784";
            when 783 => reg3_string <= " 783";
            when 782 => reg3_string <= " 782";
            when 781 => reg3_string <= " 781";
            when 780 => reg3_string <= " 780";
            when 779 => reg3_string <= " 779";
            when 778 => reg3_string <= " 778";
            when 777 => reg3_string <= " 777";
            when 776 => reg3_string <= " 776";
            when 775 => reg3_string <= " 775";
            when 774 => reg3_string <= " 774";
            when 773 => reg3_string <= " 773";
            when 772 => reg3_string <= " 772";
            when 771 => reg3_string <= " 771";
            when 770 => reg3_string <= " 770";
            when 769 => reg3_string <= " 769";
            when 768 => reg3_string <= " 768";
            when 767 => reg3_string <= " 767";
            when 766 => reg3_string <= " 766";
            when 765 => reg3_string <= " 765";
            when 764 => reg3_string <= " 764";
            when 763 => reg3_string <= " 763";
            when 762 => reg3_string <= " 762";
            when 761 => reg3_string <= " 761";
            when 760 => reg3_string <= " 760";
            when 759 => reg3_string <= " 759";
            when 758 => reg3_string <= " 758";
            when 757 => reg3_string <= " 757";
            when 756 => reg3_string <= " 756";
            when 755 => reg3_string <= " 755";
            when 754 => reg3_string <= " 754";
            when 753 => reg3_string <= " 753";
            when 752 => reg3_string <= " 752";
            when 751 => reg3_string <= " 751";
            when 750 => reg3_string <= " 750";
            when 749 => reg3_string <= " 749";
            when 748 => reg3_string <= " 748";
            when 747 => reg3_string <= " 747";
            when 746 => reg3_string <= " 746";
            when 745 => reg3_string <= " 745";
            when 744 => reg3_string <= " 744";
            when 743 => reg3_string <= " 743";
            when 742 => reg3_string <= " 742";
            when 741 => reg3_string <= " 741";
            when 740 => reg3_string <= " 740";
            when 739 => reg3_string <= " 739";
            when 738 => reg3_string <= " 738";
            when 737 => reg3_string <= " 737";
            when 736 => reg3_string <= " 736";
            when 735 => reg3_string <= " 735";
            when 734 => reg3_string <= " 734";
            when 733 => reg3_string <= " 733";
            when 732 => reg3_string <= " 732";
            when 731 => reg3_string <= " 731";
            when 730 => reg3_string <= " 730";
            when 729 => reg3_string <= " 729";
            when 728 => reg3_string <= " 728";
            when 727 => reg3_string <= " 727";
            when 726 => reg3_string <= " 726";
            when 725 => reg3_string <= " 725";
            when 724 => reg3_string <= " 724";
            when 723 => reg3_string <= " 723";
            when 722 => reg3_string <= " 722";
            when 721 => reg3_string <= " 721";
            when 720 => reg3_string <= " 720";
            when 719 => reg3_string <= " 719";
            when 718 => reg3_string <= " 718";
            when 717 => reg3_string <= " 717";
            when 716 => reg3_string <= " 716";
            when 715 => reg3_string <= " 715";
            when 714 => reg3_string <= " 714";
            when 713 => reg3_string <= " 713";
            when 712 => reg3_string <= " 712";
            when 711 => reg3_string <= " 711";
            when 710 => reg3_string <= " 710";
            when 709 => reg3_string <= " 709";
            when 708 => reg3_string <= " 708";
            when 707 => reg3_string <= " 707";
            when 706 => reg3_string <= " 706";
            when 705 => reg3_string <= " 705";
            when 704 => reg3_string <= " 704";
            when 703 => reg3_string <= " 703";
            when 702 => reg3_string <= " 702";
            when 701 => reg3_string <= " 701";
            when 700 => reg3_string <= " 700";
            when 699 => reg3_string <= " 699";
            when 698 => reg3_string <= " 698";
            when 697 => reg3_string <= " 697";
            when 696 => reg3_string <= " 696";
            when 695 => reg3_string <= " 695";
            when 694 => reg3_string <= " 694";
            when 693 => reg3_string <= " 693";
            when 692 => reg3_string <= " 692";
            when 691 => reg3_string <= " 691";
            when 690 => reg3_string <= " 690";
            when 689 => reg3_string <= " 689";
            when 688 => reg3_string <= " 688";
            when 687 => reg3_string <= " 687";
            when 686 => reg3_string <= " 686";
            when 685 => reg3_string <= " 685";
            when 684 => reg3_string <= " 684";
            when 683 => reg3_string <= " 683";
            when 682 => reg3_string <= " 682";
            when 681 => reg3_string <= " 681";
            when 680 => reg3_string <= " 680";
            when 679 => reg3_string <= " 679";
            when 678 => reg3_string <= " 678";
            when 677 => reg3_string <= " 677";
            when 676 => reg3_string <= " 676";
            when 675 => reg3_string <= " 675";
            when 674 => reg3_string <= " 674";
            when 673 => reg3_string <= " 673";
            when 672 => reg3_string <= " 672";
            when 671 => reg3_string <= " 671";
            when 670 => reg3_string <= " 670";
            when 669 => reg3_string <= " 669";
            when 668 => reg3_string <= " 668";
            when 667 => reg3_string <= " 667";
            when 666 => reg3_string <= " 666";
            when 665 => reg3_string <= " 665";
            when 664 => reg3_string <= " 664";
            when 663 => reg3_string <= " 663";
            when 662 => reg3_string <= " 662";
            when 661 => reg3_string <= " 661";
            when 660 => reg3_string <= " 660";
            when 659 => reg3_string <= " 659";
            when 658 => reg3_string <= " 658";
            when 657 => reg3_string <= " 657";
            when 656 => reg3_string <= " 656";
            when 655 => reg3_string <= " 655";
            when 654 => reg3_string <= " 654";
            when 653 => reg3_string <= " 653";
            when 652 => reg3_string <= " 652";
            when 651 => reg3_string <= " 651";
            when 650 => reg3_string <= " 650";
            when 649 => reg3_string <= " 649";
            when 648 => reg3_string <= " 648";
            when 647 => reg3_string <= " 647";
            when 646 => reg3_string <= " 646";
            when 645 => reg3_string <= " 645";
            when 644 => reg3_string <= " 644";
            when 643 => reg3_string <= " 643";
            when 642 => reg3_string <= " 642";
            when 641 => reg3_string <= " 641";
            when 640 => reg3_string <= " 640";
            when 639 => reg3_string <= " 639";
            when 638 => reg3_string <= " 638";
            when 637 => reg3_string <= " 637";
            when 636 => reg3_string <= " 636";
            when 635 => reg3_string <= " 635";
            when 634 => reg3_string <= " 634";
            when 633 => reg3_string <= " 633";
            when 632 => reg3_string <= " 632";
            when 631 => reg3_string <= " 631";
            when 630 => reg3_string <= " 630";
            when 629 => reg3_string <= " 629";
            when 628 => reg3_string <= " 628";
            when 627 => reg3_string <= " 627";
            when 626 => reg3_string <= " 626";
            when 625 => reg3_string <= " 625";
            when 624 => reg3_string <= " 624";
            when 623 => reg3_string <= " 623";
            when 622 => reg3_string <= " 622";
            when 621 => reg3_string <= " 621";
            when 620 => reg3_string <= " 620";
            when 619 => reg3_string <= " 619";
            when 618 => reg3_string <= " 618";
            when 617 => reg3_string <= " 617";
            when 616 => reg3_string <= " 616";
            when 615 => reg3_string <= " 615";
            when 614 => reg3_string <= " 614";
            when 613 => reg3_string <= " 613";
            when 612 => reg3_string <= " 612";
            when 611 => reg3_string <= " 611";
            when 610 => reg3_string <= " 610";
            when 609 => reg3_string <= " 609";
            when 608 => reg3_string <= " 608";
            when 607 => reg3_string <= " 607";
            when 606 => reg3_string <= " 606";
            when 605 => reg3_string <= " 605";
            when 604 => reg3_string <= " 604";
            when 603 => reg3_string <= " 603";
            when 602 => reg3_string <= " 602";
            when 601 => reg3_string <= " 601";
            when 600 => reg3_string <= " 600";
            when 599 => reg3_string <= " 599";
            when 598 => reg3_string <= " 598";
            when 597 => reg3_string <= " 597";
            when 596 => reg3_string <= " 596";
            when 595 => reg3_string <= " 595";
            when 594 => reg3_string <= " 594";
            when 593 => reg3_string <= " 593";
            when 592 => reg3_string <= " 592";
            when 591 => reg3_string <= " 591";
            when 590 => reg3_string <= " 590";
            when 589 => reg3_string <= " 589";
            when 588 => reg3_string <= " 588";
            when 587 => reg3_string <= " 587";
            when 586 => reg3_string <= " 586";
            when 585 => reg3_string <= " 585";
            when 584 => reg3_string <= " 584";
            when 583 => reg3_string <= " 583";
            when 582 => reg3_string <= " 582";
            when 581 => reg3_string <= " 581";
            when 580 => reg3_string <= " 580";
            when 579 => reg3_string <= " 579";
            when 578 => reg3_string <= " 578";
            when 577 => reg3_string <= " 577";
            when 576 => reg3_string <= " 576";
            when 575 => reg3_string <= " 575";
            when 574 => reg3_string <= " 574";
            when 573 => reg3_string <= " 573";
            when 572 => reg3_string <= " 572";
            when 571 => reg3_string <= " 571";
            when 570 => reg3_string <= " 570";
            when 569 => reg3_string <= " 569";
            when 568 => reg3_string <= " 568";
            when 567 => reg3_string <= " 567";
            when 566 => reg3_string <= " 566";
            when 565 => reg3_string <= " 565";
            when 564 => reg3_string <= " 564";
            when 563 => reg3_string <= " 563";
            when 562 => reg3_string <= " 562";
            when 561 => reg3_string <= " 561";
            when 560 => reg3_string <= " 560";
            when 559 => reg3_string <= " 559";
            when 558 => reg3_string <= " 558";
            when 557 => reg3_string <= " 557";
            when 556 => reg3_string <= " 556";
            when 555 => reg3_string <= " 555";
            when 554 => reg3_string <= " 554";
            when 553 => reg3_string <= " 553";
            when 552 => reg3_string <= " 552";
            when 551 => reg3_string <= " 551";
            when 550 => reg3_string <= " 550";
            when 549 => reg3_string <= " 549";
            when 548 => reg3_string <= " 548";
            when 547 => reg3_string <= " 547";
            when 546 => reg3_string <= " 546";
            when 545 => reg3_string <= " 545";
            when 544 => reg3_string <= " 544";
            when 543 => reg3_string <= " 543";
            when 542 => reg3_string <= " 542";
            when 541 => reg3_string <= " 541";
            when 540 => reg3_string <= " 540";
            when 539 => reg3_string <= " 539";
            when 538 => reg3_string <= " 538";
            when 537 => reg3_string <= " 537";
            when 536 => reg3_string <= " 536";
            when 535 => reg3_string <= " 535";
            when 534 => reg3_string <= " 534";
            when 533 => reg3_string <= " 533";
            when 532 => reg3_string <= " 532";
            when 531 => reg3_string <= " 531";
            when 530 => reg3_string <= " 530";
            when 529 => reg3_string <= " 529";
            when 528 => reg3_string <= " 528";
            when 527 => reg3_string <= " 527";
            when 526 => reg3_string <= " 526";
            when 525 => reg3_string <= " 525";
            when 524 => reg3_string <= " 524";
            when 523 => reg3_string <= " 523";
            when 522 => reg3_string <= " 522";
            when 521 => reg3_string <= " 521";
            when 520 => reg3_string <= " 520";
            when 519 => reg3_string <= " 519";
            when 518 => reg3_string <= " 518";
            when 517 => reg3_string <= " 517";
            when 516 => reg3_string <= " 516";
            when 515 => reg3_string <= " 515";
            when 514 => reg3_string <= " 514";
            when 513 => reg3_string <= " 513";
            when 512 => reg3_string <= " 512";
            when 511 => reg3_string <= " 511";
            when 510 => reg3_string <= " 510";
            when 509 => reg3_string <= " 509";
            when 508 => reg3_string <= " 508";
            when 507 => reg3_string <= " 507";
            when 506 => reg3_string <= " 506";
            when 505 => reg3_string <= " 505";
            when 504 => reg3_string <= " 504";
            when 503 => reg3_string <= " 503";
            when 502 => reg3_string <= " 502";
            when 501 => reg3_string <= " 501";
            when 500 => reg3_string <= " 500";
            when 499 => reg3_string <= " 499";
            when 498 => reg3_string <= " 498";
            when 497 => reg3_string <= " 497";
            when 496 => reg3_string <= " 496";
            when 495 => reg3_string <= " 495";
            when 494 => reg3_string <= " 494";
            when 493 => reg3_string <= " 493";
            when 492 => reg3_string <= " 492";
            when 491 => reg3_string <= " 491";
            when 490 => reg3_string <= " 490";
            when 489 => reg3_string <= " 489";
            when 488 => reg3_string <= " 488";
            when 487 => reg3_string <= " 487";
            when 486 => reg3_string <= " 486";
            when 485 => reg3_string <= " 485";
            when 484 => reg3_string <= " 484";
            when 483 => reg3_string <= " 483";
            when 482 => reg3_string <= " 482";
            when 481 => reg3_string <= " 481";
            when 480 => reg3_string <= " 480";
            when 479 => reg3_string <= " 479";
            when 478 => reg3_string <= " 478";
            when 477 => reg3_string <= " 477";
            when 476 => reg3_string <= " 476";
            when 475 => reg3_string <= " 475";
            when 474 => reg3_string <= " 474";
            when 473 => reg3_string <= " 473";
            when 472 => reg3_string <= " 472";
            when 471 => reg3_string <= " 471";
            when 470 => reg3_string <= " 470";
            when 469 => reg3_string <= " 469";
            when 468 => reg3_string <= " 468";
            when 467 => reg3_string <= " 467";
            when 466 => reg3_string <= " 466";
            when 465 => reg3_string <= " 465";
            when 464 => reg3_string <= " 464";
            when 463 => reg3_string <= " 463";
            when 462 => reg3_string <= " 462";
            when 461 => reg3_string <= " 461";
            when 460 => reg3_string <= " 460";
            when 459 => reg3_string <= " 459";
            when 458 => reg3_string <= " 458";
            when 457 => reg3_string <= " 457";
            when 456 => reg3_string <= " 456";
            when 455 => reg3_string <= " 455";
            when 454 => reg3_string <= " 454";
            when 453 => reg3_string <= " 453";
            when 452 => reg3_string <= " 452";
            when 451 => reg3_string <= " 451";
            when 450 => reg3_string <= " 450";
            when 449 => reg3_string <= " 449";
            when 448 => reg3_string <= " 448";
            when 447 => reg3_string <= " 447";
            when 446 => reg3_string <= " 446";
            when 445 => reg3_string <= " 445";
            when 444 => reg3_string <= " 444";
            when 443 => reg3_string <= " 443";
            when 442 => reg3_string <= " 442";
            when 441 => reg3_string <= " 441";
            when 440 => reg3_string <= " 440";
            when 439 => reg3_string <= " 439";
            when 438 => reg3_string <= " 438";
            when 437 => reg3_string <= " 437";
            when 436 => reg3_string <= " 436";
            when 435 => reg3_string <= " 435";
            when 434 => reg3_string <= " 434";
            when 433 => reg3_string <= " 433";
            when 432 => reg3_string <= " 432";
            when 431 => reg3_string <= " 431";
            when 430 => reg3_string <= " 430";
            when 429 => reg3_string <= " 429";
            when 428 => reg3_string <= " 428";
            when 427 => reg3_string <= " 427";
            when 426 => reg3_string <= " 426";
            when 425 => reg3_string <= " 425";
            when 424 => reg3_string <= " 424";
            when 423 => reg3_string <= " 423";
            when 422 => reg3_string <= " 422";
            when 421 => reg3_string <= " 421";
            when 420 => reg3_string <= " 420";
            when 419 => reg3_string <= " 419";
            when 418 => reg3_string <= " 418";
            when 417 => reg3_string <= " 417";
            when 416 => reg3_string <= " 416";
            when 415 => reg3_string <= " 415";
            when 414 => reg3_string <= " 414";
            when 413 => reg3_string <= " 413";
            when 412 => reg3_string <= " 412";
            when 411 => reg3_string <= " 411";
            when 410 => reg3_string <= " 410";
            when 409 => reg3_string <= " 409";
            when 408 => reg3_string <= " 408";
            when 407 => reg3_string <= " 407";
            when 406 => reg3_string <= " 406";
            when 405 => reg3_string <= " 405";
            when 404 => reg3_string <= " 404";
            when 403 => reg3_string <= " 403";
            when 402 => reg3_string <= " 402";
            when 401 => reg3_string <= " 401";
            when 400 => reg3_string <= " 400";
            when 399 => reg3_string <= " 399";
            when 398 => reg3_string <= " 398";
            when 397 => reg3_string <= " 397";
            when 396 => reg3_string <= " 396";
            when 395 => reg3_string <= " 395";
            when 394 => reg3_string <= " 394";
            when 393 => reg3_string <= " 393";
            when 392 => reg3_string <= " 392";
            when 391 => reg3_string <= " 391";
            when 390 => reg3_string <= " 390";
            when 389 => reg3_string <= " 389";
            when 388 => reg3_string <= " 388";
            when 387 => reg3_string <= " 387";
            when 386 => reg3_string <= " 386";
            when 385 => reg3_string <= " 385";
            when 384 => reg3_string <= " 384";
            when 383 => reg3_string <= " 383";
            when 382 => reg3_string <= " 382";
            when 381 => reg3_string <= " 381";
            when 380 => reg3_string <= " 380";
            when 379 => reg3_string <= " 379";
            when 378 => reg3_string <= " 378";
            when 377 => reg3_string <= " 377";
            when 376 => reg3_string <= " 376";
            when 375 => reg3_string <= " 375";
            when 374 => reg3_string <= " 374";
            when 373 => reg3_string <= " 373";
            when 372 => reg3_string <= " 372";
            when 371 => reg3_string <= " 371";
            when 370 => reg3_string <= " 370";
            when 369 => reg3_string <= " 369";
            when 368 => reg3_string <= " 368";
            when 367 => reg3_string <= " 367";
            when 366 => reg3_string <= " 366";
            when 365 => reg3_string <= " 365";
            when 364 => reg3_string <= " 364";
            when 363 => reg3_string <= " 363";
            when 362 => reg3_string <= " 362";
            when 361 => reg3_string <= " 361";
            when 360 => reg3_string <= " 360";
            when 359 => reg3_string <= " 359";
            when 358 => reg3_string <= " 358";
            when 357 => reg3_string <= " 357";
            when 356 => reg3_string <= " 356";
            when 355 => reg3_string <= " 355";
            when 354 => reg3_string <= " 354";
            when 353 => reg3_string <= " 353";
            when 352 => reg3_string <= " 352";
            when 351 => reg3_string <= " 351";
            when 350 => reg3_string <= " 350";
            when 349 => reg3_string <= " 349";
            when 348 => reg3_string <= " 348";
            when 347 => reg3_string <= " 347";
            when 346 => reg3_string <= " 346";
            when 345 => reg3_string <= " 345";
            when 344 => reg3_string <= " 344";
            when 343 => reg3_string <= " 343";
            when 342 => reg3_string <= " 342";
            when 341 => reg3_string <= " 341";
            when 340 => reg3_string <= " 340";
            when 339 => reg3_string <= " 339";
            when 338 => reg3_string <= " 338";
            when 337 => reg3_string <= " 337";
            when 336 => reg3_string <= " 336";
            when 335 => reg3_string <= " 335";
            when 334 => reg3_string <= " 334";
            when 333 => reg3_string <= " 333";
            when 332 => reg3_string <= " 332";
            when 331 => reg3_string <= " 331";
            when 330 => reg3_string <= " 330";
            when 329 => reg3_string <= " 329";
            when 328 => reg3_string <= " 328";
            when 327 => reg3_string <= " 327";
            when 326 => reg3_string <= " 326";
            when 325 => reg3_string <= " 325";
            when 324 => reg3_string <= " 324";
            when 323 => reg3_string <= " 323";
            when 322 => reg3_string <= " 322";
            when 321 => reg3_string <= " 321";
            when 320 => reg3_string <= " 320";
            when 319 => reg3_string <= " 319";
            when 318 => reg3_string <= " 318";
            when 317 => reg3_string <= " 317";
            when 316 => reg3_string <= " 316";
            when 315 => reg3_string <= " 315";
            when 314 => reg3_string <= " 314";
            when 313 => reg3_string <= " 313";
            when 312 => reg3_string <= " 312";
            when 311 => reg3_string <= " 311";
            when 310 => reg3_string <= " 310";
            when 309 => reg3_string <= " 309";
            when 308 => reg3_string <= " 308";
            when 307 => reg3_string <= " 307";
            when 306 => reg3_string <= " 306";
            when 305 => reg3_string <= " 305";
            when 304 => reg3_string <= " 304";
            when 303 => reg3_string <= " 303";
            when 302 => reg3_string <= " 302";
            when 301 => reg3_string <= " 301";
            when 300 => reg3_string <= " 300";
            when 299 => reg3_string <= " 299";
            when 298 => reg3_string <= " 298";
            when 297 => reg3_string <= " 297";
            when 296 => reg3_string <= " 296";
            when 295 => reg3_string <= " 295";
            when 294 => reg3_string <= " 294";
            when 293 => reg3_string <= " 293";
            when 292 => reg3_string <= " 292";
            when 291 => reg3_string <= " 291";
            when 290 => reg3_string <= " 290";
            when 289 => reg3_string <= " 289";
            when 288 => reg3_string <= " 288";
            when 287 => reg3_string <= " 287";
            when 286 => reg3_string <= " 286";
            when 285 => reg3_string <= " 285";
            when 284 => reg3_string <= " 284";
            when 283 => reg3_string <= " 283";
            when 282 => reg3_string <= " 282";
            when 281 => reg3_string <= " 281";
            when 280 => reg3_string <= " 280";
            when 279 => reg3_string <= " 279";
            when 278 => reg3_string <= " 278";
            when 277 => reg3_string <= " 277";
            when 276 => reg3_string <= " 276";
            when 275 => reg3_string <= " 275";
            when 274 => reg3_string <= " 274";
            when 273 => reg3_string <= " 273";
            when 272 => reg3_string <= " 272";
            when 271 => reg3_string <= " 271";
            when 270 => reg3_string <= " 270";
            when 269 => reg3_string <= " 269";
            when 268 => reg3_string <= " 268";
            when 267 => reg3_string <= " 267";
            when 266 => reg3_string <= " 266";
            when 265 => reg3_string <= " 265";
            when 264 => reg3_string <= " 264";
            when 263 => reg3_string <= " 263";
            when 262 => reg3_string <= " 262";
            when 261 => reg3_string <= " 261";
            when 260 => reg3_string <= " 260";
            when 259 => reg3_string <= " 259";
            when 258 => reg3_string <= " 258";
            when 257 => reg3_string <= " 257";
            when 256 => reg3_string <= " 256";
            when 255 => reg3_string <= " 255";
            when 254 => reg3_string <= " 254";
            when 253 => reg3_string <= " 253";
            when 252 => reg3_string <= " 252";
            when 251 => reg3_string <= " 251";
            when 250 => reg3_string <= " 250";
            when 249 => reg3_string <= " 249";
            when 248 => reg3_string <= " 248";
            when 247 => reg3_string <= " 247";
            when 246 => reg3_string <= " 246";
            when 245 => reg3_string <= " 245";
            when 244 => reg3_string <= " 244";
            when 243 => reg3_string <= " 243";
            when 242 => reg3_string <= " 242";
            when 241 => reg3_string <= " 241";
            when 240 => reg3_string <= " 240";
            when 239 => reg3_string <= " 239";
            when 238 => reg3_string <= " 238";
            when 237 => reg3_string <= " 237";
            when 236 => reg3_string <= " 236";
            when 235 => reg3_string <= " 235";
            when 234 => reg3_string <= " 234";
            when 233 => reg3_string <= " 233";
            when 232 => reg3_string <= " 232";
            when 231 => reg3_string <= " 231";
            when 230 => reg3_string <= " 230";
            when 229 => reg3_string <= " 229";
            when 228 => reg3_string <= " 228";
            when 227 => reg3_string <= " 227";
            when 226 => reg3_string <= " 226";
            when 225 => reg3_string <= " 225";
            when 224 => reg3_string <= " 224";
            when 223 => reg3_string <= " 223";
            when 222 => reg3_string <= " 222";
            when 221 => reg3_string <= " 221";
            when 220 => reg3_string <= " 220";
            when 219 => reg3_string <= " 219";
            when 218 => reg3_string <= " 218";
            when 217 => reg3_string <= " 217";
            when 216 => reg3_string <= " 216";
            when 215 => reg3_string <= " 215";
            when 214 => reg3_string <= " 214";
            when 213 => reg3_string <= " 213";
            when 212 => reg3_string <= " 212";
            when 211 => reg3_string <= " 211";
            when 210 => reg3_string <= " 210";
            when 209 => reg3_string <= " 209";
            when 208 => reg3_string <= " 208";
            when 207 => reg3_string <= " 207";
            when 206 => reg3_string <= " 206";
            when 205 => reg3_string <= " 205";
            when 204 => reg3_string <= " 204";
            when 203 => reg3_string <= " 203";
            when 202 => reg3_string <= " 202";
            when 201 => reg3_string <= " 201";
            when 200 => reg3_string <= " 200";
            when 199 => reg3_string <= " 199";
            when 198 => reg3_string <= " 198";
            when 197 => reg3_string <= " 197";
            when 196 => reg3_string <= " 196";
            when 195 => reg3_string <= " 195";
            when 194 => reg3_string <= " 194";
            when 193 => reg3_string <= " 193";
            when 192 => reg3_string <= " 192";
            when 191 => reg3_string <= " 191";
            when 190 => reg3_string <= " 190";
            when 189 => reg3_string <= " 189";
            when 188 => reg3_string <= " 188";
            when 187 => reg3_string <= " 187";
            when 186 => reg3_string <= " 186";
            when 185 => reg3_string <= " 185";
            when 184 => reg3_string <= " 184";
            when 183 => reg3_string <= " 183";
            when 182 => reg3_string <= " 182";
            when 181 => reg3_string <= " 181";
            when 180 => reg3_string <= " 180";
            when 179 => reg3_string <= " 179";
            when 178 => reg3_string <= " 178";
            when 177 => reg3_string <= " 177";
            when 176 => reg3_string <= " 176";
            when 175 => reg3_string <= " 175";
            when 174 => reg3_string <= " 174";
            when 173 => reg3_string <= " 173";
            when 172 => reg3_string <= " 172";
            when 171 => reg3_string <= " 171";
            when 170 => reg3_string <= " 170";
            when 169 => reg3_string <= " 169";
            when 168 => reg3_string <= " 168";
            when 167 => reg3_string <= " 167";
            when 166 => reg3_string <= " 166";
            when 165 => reg3_string <= " 165";
            when 164 => reg3_string <= " 164";
            when 163 => reg3_string <= " 163";
            when 162 => reg3_string <= " 162";
            when 161 => reg3_string <= " 161";
            when 160 => reg3_string <= " 160";
            when 159 => reg3_string <= " 159";
            when 158 => reg3_string <= " 158";
            when 157 => reg3_string <= " 157";
            when 156 => reg3_string <= " 156";
            when 155 => reg3_string <= " 155";
            when 154 => reg3_string <= " 154";
            when 153 => reg3_string <= " 153";
            when 152 => reg3_string <= " 152";
            when 151 => reg3_string <= " 151";
            when 150 => reg3_string <= " 150";
            when 149 => reg3_string <= " 149";
            when 148 => reg3_string <= " 148";
            when 147 => reg3_string <= " 147";
            when 146 => reg3_string <= " 146";
            when 145 => reg3_string <= " 145";
            when 144 => reg3_string <= " 144";
            when 143 => reg3_string <= " 143";
            when 142 => reg3_string <= " 142";
            when 141 => reg3_string <= " 141";
            when 140 => reg3_string <= " 140";
            when 139 => reg3_string <= " 139";
            when 138 => reg3_string <= " 138";
            when 137 => reg3_string <= " 137";
            when 136 => reg3_string <= " 136";
            when 135 => reg3_string <= " 135";
            when 134 => reg3_string <= " 134";
            when 133 => reg3_string <= " 133";
            when 132 => reg3_string <= " 132";
            when 131 => reg3_string <= " 131";
            when 130 => reg3_string <= " 130";
            when 129 => reg3_string <= " 129";
            when 128 => reg3_string <= " 128";
            when 127 => reg3_string <= " 127";
            when 126 => reg3_string <= " 126";
            when 125 => reg3_string <= " 125";
            when 124 => reg3_string <= " 124";
            when 123 => reg3_string <= " 123";
            when 122 => reg3_string <= " 122";
            when 121 => reg3_string <= " 121";
            when 120 => reg3_string <= " 120";
            when 119 => reg3_string <= " 119";
            when 118 => reg3_string <= " 118";
            when 117 => reg3_string <= " 117";
            when 116 => reg3_string <= " 116";
            when 115 => reg3_string <= " 115";
            when 114 => reg3_string <= " 114";
            when 113 => reg3_string <= " 113";
            when 112 => reg3_string <= " 112";
            when 111 => reg3_string <= " 111";
            when 110 => reg3_string <= " 110";
            when 109 => reg3_string <= " 109";
            when 108 => reg3_string <= " 108";
            when 107 => reg3_string <= " 107";                                                                                        
            when 106 => reg3_string <= " 106";                                                                                        
            when 105 => reg3_string <= " 105";                                                                                        
            when 104 => reg3_string <= " 104";                                                                                        
            when 103 => reg3_string <= " 103";                                                                                        
            when 102 => reg3_string <= " 102";                                                                                        
            when 101 => reg3_string <= " 101";                                                                                        
            when 100 => reg3_string <= " 100";                                                                                        
            when 99 => reg3_string <= "  99";                                                                                         
            when 98 => reg3_string <= "  98";                                                                                         
            when 97 => reg3_string <= "  97";                                                                                         
            when 96 => reg3_string <= "  96";                                                                                         
            when 95 => reg3_string <= "  95";                                                                                         
            when 94 => reg3_string <= "  94";                                                                                         
            when 93 => reg3_string <= "  93";                                                                                         
            when 92 => reg3_string <= "  92";                                                                                         
            when 91 => reg3_string <= "  91";                                                                                         
            when 90 => reg3_string <= "  90";                                                                                         
            when 89 => reg3_string <= "  89";                                                                                         
            when 88 => reg3_string <= "  88";                                                                                         
            when 87 => reg3_string <= "  87";                                                                                         
            when 86 => reg3_string <= "  86";                                                                                         
            when 85 => reg3_string <= "  85";                                                                                         
            when 84 => reg3_string <= "  84";                                                                                         
            when 83 => reg3_string <= "  83";                                                                                         
            when 82 => reg3_string <= "  82";                                                                                         
            when 81 => reg3_string <= "  81";                                                                                         
            when 80 => reg3_string <= "  80";                                                                                         
            when 79 => reg3_string <= "  79";                                                                                         
            when 78 => reg3_string <= "  78";                                                                                         
            when 77 => reg3_string <= "  77";  
            when 76 => reg3_string <= "  76";                                                                                         
            when 75 => reg3_string <= "  75";                                                                                         
            when 74 => reg3_string <= "  74";                                                                                         
            when 73 => reg3_string <= "  73";                                                                                         
            when 72 => reg3_string <= "  72";                                                                                         
            when 71 => reg3_string <= "  71";                                                                                         
            when 70 => reg3_string <= "  70";                                                                                         
            when 69 => reg3_string <= "  69";                                                                                         
            when 68 => reg3_string <= "  68";                                                                                         
            when 67 => reg3_string <= "  67";                                                                                         
            when 66 => reg3_string <= "  66";                                                                                         
            when 65 => reg3_string <= "  65";                                                                                         
            when 64 => reg3_string <= "  64";                                                                                         
            when 63 => reg3_string <= "  63";                                                                                         
            when 62 => reg3_string <= "  62";                                                                                         
            when 61 => reg3_string <= "  61";                                                                                         
            when 60 => reg3_string <= "  60";                                                                                         
            when 59 => reg3_string <= "  59";                                                                                         
            when 58 => reg3_string <= "  58";                                                                                         
            when 57 => reg3_string <= "  57";                                                                                         
            when 56 => reg3_string <= "  56";                                                                                         
            when 55 => reg3_string <= "  55";                                                                                         
            when 54 => reg3_string <= "  54";                                                                                         
            when 53 => reg3_string <= "  53";                                                                                         
            when 52 => reg3_string <= "  52";                                                                                         
            when 51 => reg3_string <= "  51";                                                                                         
            when 50 => reg3_string <= "  50";                                                                                         
            when 49 => reg3_string <= "  49";                                                                                         
            when 48 => reg3_string <= "  48";                                                                                         
            when 47 => reg3_string <= "  47";
            when 46 => reg3_string <= "  46";                                                                                         
            when 45 => reg3_string <= "  45";                                                                                         
            when 44 => reg3_string <= "  44";                                                                                         
            when 43 => reg3_string <= "  43";                                                                                         
            when 42 => reg3_string <= "  42";                                                                                         
            when 41 => reg3_string <= "  41";                                                                                         
            when 40 => reg3_string <= "  40";                                                                                         
            when 39 => reg3_string <= "  39";                                                                                         
            when 38 => reg3_string <= "  38";                                                                                         
            when 37 => reg3_string <= "  37";                                                                                         
            when 36 => reg3_string <= "  36";                                                                                         
            when 35 => reg3_string <= "  35";                                                                                         
            when 34 => reg3_string <= "  34";                                                                                         
            when 33 => reg3_string <= "  33";                                                                                         
            when 32 => reg3_string <= "  32";                                                                                         
            when 31 => reg3_string <= "  31";                                                                                         
            when 30 => reg3_string <= "  30";                                                                                         
            when 29 => reg3_string <= "  29";                                                                                         
            when 28 => reg3_string <= "  28";                                                                                         
            when 27 => reg3_string <= "  27";                                                                                         
            when 26 => reg3_string <= "  26";                                                                                         
            when 25 => reg3_string <= "  25";                                                                                         
            when 24 => reg3_string <= "  24";                                                                                         
            when 23 => reg3_string <= "  23";
            when 22 => reg3_string <= "  22";                                                                                         
            when 21 => reg3_string <= "  21";                                                                                         
            when 20 => reg3_string <= "  20";                                                                                         
            when 19 => reg3_string <= "  19";                                                                                         
            when 18 => reg3_string <= "  18";                                                                                         
            when 17 => reg3_string <= "  17";                                                                                         
            when 16 => reg3_string <= "  16";                                                                                         
            when 15 => reg3_string <= "  15";                                                                                         
            when 14 => reg3_string <= "  14";                                                                                         
            when 13 => reg3_string <= "  13";                                                                                         
            when 12 => reg3_string <= "  12";                                                                                         
            when 11 => reg3_string <= "  11";                                                                                         
            when 10 => reg3_string <= "  10";                                                                                         
            when 9  => reg3_string <= "   9";                                                                                          
            when 8  => reg3_string <= "   8";                                                                                          
            when 7  => reg3_string <= "   7";                                                                                          
            when 6  => reg3_string <= "   6";                                                                                          
            when 5  => reg3_string <= "   5";                                                                                          
            when 4  => reg3_string <= "   4";                                                                                          
            when 3  => reg3_string <= "   3";                                                                                          
            when 2  => reg3_string <= "   2";                                                                                          
            when 1  => reg3_string <= "   1";                                                                                          
            when 0  => reg3_string <= "   0";
            when -1 => reg3_string <= "  -1";
            when -2 => reg3_string <= "  -2";
            when -3 => reg3_string <= "  -3";
            when -4 => reg3_string <= "  -4";
            when -5 => reg3_string <= "  -5";
            when -6 => reg3_string <= "  -6";
            when -7 => reg3_string <= "  -7";
            when -8 => reg3_string <= "  -8";
            when -9 => reg3_string <= "  -9";
            when -10 => reg3_string <= " -10";
            when -11 => reg3_string <= " -11";
            when -12 => reg3_string <= " -12";
            when -13 => reg3_string <= " -13";
            when -14 => reg3_string <= " -14";
            when -15 => reg3_string <= " -15";
            when -16 => reg3_string <= " -16";
            when -17 => reg3_string <= " -17";
            when -18 => reg3_string <= " -18";
            when -19 => reg3_string <= " -19";
            when -20 => reg3_string <= " -20";
            when -21 => reg3_string <= " -21";
            when -22 => reg3_string <= " -22";
            when -23 => reg3_string <= " -23";
            when -24 => reg3_string <= " -24";
            when -25 => reg3_string <= " -25";
            when -26 => reg3_string <= " -26";
            when -27 => reg3_string <= " -27";
            when -28 => reg3_string <= " -28";
            when -29 => reg3_string <= " -29";
            when -30 => reg3_string <= " -30";
            when -31 => reg3_string <= " -31";
            when -32 => reg3_string <= " -32";
            when -33 => reg3_string <= " -33";
            when -34 => reg3_string <= " -34";
            when -35 => reg3_string <= " -35";
            when -36 => reg3_string <= " -36";
            when -37 => reg3_string <= " -37";
            when -38 => reg3_string <= " -38";
            when -39 => reg3_string <= " -39";
            when -40 => reg3_string <= " -40";
            when -41 => reg3_string <= " -41";
            when -42 => reg3_string <= " -42";
            when -43 => reg3_string <= " -43";
            when -44 => reg3_string <= " -44";
            when -45 => reg3_string <= " -45";
            when -46 => reg3_string <= " -46";
            when -47 => reg3_string <= " -47";
            when -48 => reg3_string <= " -48";
            when -49 => reg3_string <= " -49";
            when -50 => reg3_string <= " -50";
            when -51 => reg3_string <= " -51";
            when -52 => reg3_string <= " -52";
            when -53 => reg3_string <= " -53";
            when -54 => reg3_string <= " -54";
            when -55 => reg3_string <= " -55";
            when -56 => reg3_string <= " -56";
            when -57 => reg3_string <= " -57";
            when -58 => reg3_string <= " -58";
            when -59 => reg3_string <= " -59";
            when -60 => reg3_string <= " -60";
            when -61 => reg3_string <= " -61";
            when -62 => reg3_string <= " -62";
            when -63 => reg3_string <= " -63";
            when -64 => reg3_string <= " -64";
            when -65 => reg3_string <= " -65";
            when -66 => reg3_string <= " -66";
            when -67 => reg3_string <= " -67";
            when -68 => reg3_string <= " -68";
            when -69 => reg3_string <= " -69";
            when -70 => reg3_string <= " -70";
            when -71 => reg3_string <= " -71";
            when -72 => reg3_string <= " -72";
            when -73 => reg3_string <= " -73";
            when -74 => reg3_string <= " -74";
            when -75 => reg3_string <= " -75";
            when -76 => reg3_string <= " -76";
            when -77 => reg3_string <= " -77";
            when -78 => reg3_string <= " -78";
            when -79 => reg3_string <= " -79";
            when -80 => reg3_string <= " -80";
            when -81 => reg3_string <= " -81";
            when -82 => reg3_string <= " -82";
            when -83 => reg3_string <= " -83";
            when -84 => reg3_string <= " -84";
            when -85 => reg3_string <= " -85";
            when -86 => reg3_string <= " -86";
            when -87 => reg3_string <= " -87";
            when -88 => reg3_string <= " -88";
            when -89 => reg3_string <= " -89";
            when -90 => reg3_string <= " -90";
            when -91 => reg3_string <= " -91";
            when -92 => reg3_string <= " -92";
            when -93 => reg3_string <= " -93";
            when -94 => reg3_string <= " -94";
            when -95 => reg3_string <= " -95";
            when -96 => reg3_string <= " -96";
            when -97 => reg3_string <= " -97";
            when -98 => reg3_string <= " -98";
            when -99 => reg3_string <= " -99";
            when -100 => reg3_string <= "-100";
            when -101 => reg3_string <= "-101";
            when -102 => reg3_string <= "-102";
            when -103 => reg3_string <= "-103";
            when -104 => reg3_string <= "-104";
            when -105 => reg3_string <= "-105";
            when -106 => reg3_string <= "-106";
            when -107 => reg3_string <= "-107";
            when -108 => reg3_string <= "-108";
            when -109 => reg3_string <= "-109";
            when -110 => reg3_string <= "-110";
            when -111 => reg3_string <= "-111";
            when -112 => reg3_string <= "-112";
            when -113 => reg3_string <= "-113";
            when -114 => reg3_string <= "-114";
            when -115 => reg3_string <= "-115";
            when -116 => reg3_string <= "-116";
            when -117 => reg3_string <= "-117";
            when -118 => reg3_string <= "-118";
            when -119 => reg3_string <= "-119";
            when -120 => reg3_string <= "-120";
            when -121 => reg3_string <= "-121";
            when -122 => reg3_string <= "-122";
            when -123 => reg3_string <= "-123";
            when -124 => reg3_string <= "-124";
            when -125 => reg3_string <= "-125";
            when -126 => reg3_string <= "-126";
            when -127 => reg3_string <= "-127";
            when -128 => reg3_string <= "-128";
            when -129 => reg3_string <= "-129";
            when -130 => reg3_string <= "-130";
            when -131 => reg3_string <= "-131";
            when -132 => reg3_string <= "-132";
            when -133 => reg3_string <= "-133";
            when -134 => reg3_string <= "-134";
            when -135 => reg3_string <= "-135";
            when -136 => reg3_string <= "-136";
            when -137 => reg3_string <= "-137";
            when -138 => reg3_string <= "-138";
            when -139 => reg3_string <= "-139";
            when -140 => reg3_string <= "-140";
            when -141 => reg3_string <= "-141";
            when -142 => reg3_string <= "-142";
            when -143 => reg3_string <= "-143";
            when -144 => reg3_string <= "-144";
            when -145 => reg3_string <= "-145";
            when -146 => reg3_string <= "-146";
            when -147 => reg3_string <= "-147";
            when -148 => reg3_string <= "-148";
            when -149 => reg3_string <= "-149";
            when -150 => reg3_string <= "-150";
            when -151 => reg3_string <= "-151";
            when -152 => reg3_string <= "-152";
            when -153 => reg3_string <= "-153";
            when -154 => reg3_string <= "-154";
            when -155 => reg3_string <= "-155";
            when -156 => reg3_string <= "-156";
            when -157 => reg3_string <= "-157";
            when -158 => reg3_string <= "-158";
            when -159 => reg3_string <= "-159";
            when -160 => reg3_string <= "-160";
            when -161 => reg3_string <= "-161";
            when -162 => reg3_string <= "-162";
            when -163 => reg3_string <= "-163";
            when -164 => reg3_string <= "-164";
            when -165 => reg3_string <= "-165";
            when -166 => reg3_string <= "-166";
            when -167 => reg3_string <= "-167";
            when -168 => reg3_string <= "-168";
            when -169 => reg3_string <= "-169";
            when -170 => reg3_string <= "-170";
            when -171 => reg3_string <= "-171";
            when -172 => reg3_string <= "-172";
            when -173 => reg3_string <= "-173";
            when -174 => reg3_string <= "-174";
            when -175 => reg3_string <= "-175";
            when -176 => reg3_string <= "-176";
            when -177 => reg3_string <= "-177";
            when -178 => reg3_string <= "-178";
            when -179 => reg3_string <= "-179";
            when -180 => reg3_string <= "-180";
            when -181 => reg3_string <= "-181";
            when -182 => reg3_string <= "-182";
            when -183 => reg3_string <= "-183";
            when -184 => reg3_string <= "-184";
            when -185 => reg3_string <= "-185";
            when -186 => reg3_string <= "-186";
            when -187 => reg3_string <= "-187";
            when -188 => reg3_string <= "-188";
            when -189 => reg3_string <= "-189";
            when -190 => reg3_string <= "-190";
            when -191 => reg3_string <= "-191";
            when -192 => reg3_string <= "-192";
            when -193 => reg3_string <= "-193";
            when -194 => reg3_string <= "-194";
            when -195 => reg3_string <= "-195";
            when -196 => reg3_string <= "-196";
            when -197 => reg3_string <= "-197";
            when -198 => reg3_string <= "-198";
            when -199 => reg3_string <= "-199";
            when -200 => reg3_string <= "-200";
            when -201 => reg3_string <= "-201";
            when -202 => reg3_string <= "-202";
            when -203 => reg3_string <= "-203";
            when -204 => reg3_string <= "-204";
            when -205 => reg3_string <= "-205";
            when -206 => reg3_string <= "-206";
            when -207 => reg3_string <= "-207";
            when -208 => reg3_string <= "-208";
            when -209 => reg3_string <= "-209";
            when -210 => reg3_string <= "-210";
            when -211 => reg3_string <= "-211";
            when -212 => reg3_string <= "-212";
            when -213 => reg3_string <= "-213";
            when -214 => reg3_string <= "-214";
            when -215 => reg3_string <= "-215";
            when -216 => reg3_string <= "-216";
            when -217 => reg3_string <= "-217";
            when -218 => reg3_string <= "-218";
            when -219 => reg3_string <= "-219";
            when -220 => reg3_string <= "-220";
            when -221 => reg3_string <= "-221";
            when -222 => reg3_string <= "-222";
            when -223 => reg3_string <= "-223";
            when -224 => reg3_string <= "-224";
            when -225 => reg3_string <= "-225";
            when -226 => reg3_string <= "-226";
            when -227 => reg3_string <= "-227";
            when -228 => reg3_string <= "-228";
            when -229 => reg3_string <= "-229";
            when -230 => reg3_string <= "-230";
            when -231 => reg3_string <= "-231";
            when -232 => reg3_string <= "-232";
            when -233 => reg3_string <= "-233";
            when -234 => reg3_string <= "-234";
            when -235 => reg3_string <= "-235";
            when -236 => reg3_string <= "-236";
            when -237 => reg3_string <= "-237";
            when -238 => reg3_string <= "-238";
            when -239 => reg3_string <= "-239";
            when -240 => reg3_string <= "-240";
            when -241 => reg3_string <= "-241";
            when -242 => reg3_string <= "-242";
            when -243 => reg3_string <= "-243";
            when -244 => reg3_string <= "-244";
            when -245 => reg3_string <= "-245";
            when -246 => reg3_string <= "-246";
            when -247 => reg3_string <= "-247";
            when -248 => reg3_string <= "-248";
            when -249 => reg3_string <= "-249";
            when -250 => reg3_string <= "-250";
            when -251 => reg3_string <= "-251";
            when -252 => reg3_string <= "-252";
            when -253 => reg3_string <= "-253";
            when -254 => reg3_string <= "-254";
            when -255 => reg3_string <= "-255";
            when -256 => reg3_string <= "-256";
            when -257 => reg3_string <= "-257";
            when -258 => reg3_string <= "-258";
            when -259 => reg3_string <= "-259";
            when -260 => reg3_string <= "-260";
            when -261 => reg3_string <= "-261";
            when -262 => reg3_string <= "-262";
            when -263 => reg3_string <= "-263";
            when -264 => reg3_string <= "-264";
            when -265 => reg3_string <= "-265";
            when -266 => reg3_string <= "-266";
            when -267 => reg3_string <= "-267";
            when -268 => reg3_string <= "-268";
            when -269 => reg3_string <= "-269";
            when -270 => reg3_string <= "-270";
            when -271 => reg3_string <= "-271";
            when -272 => reg3_string <= "-272";
            when -273 => reg3_string <= "-273";
            when -274 => reg3_string <= "-274";
            when -275 => reg3_string <= "-275";
            when -276 => reg3_string <= "-276";
            when -277 => reg3_string <= "-277";
            when -278 => reg3_string <= "-278";
            when -279 => reg3_string <= "-279";
            when -280 => reg3_string <= "-280";
            when -281 => reg3_string <= "-281";
            when -282 => reg3_string <= "-282";
            when -283 => reg3_string <= "-283";
            when -284 => reg3_string <= "-284";
            when -285 => reg3_string <= "-285";
            when -286 => reg3_string <= "-286";
            when -287 => reg3_string <= "-287";
            when -288 => reg3_string <= "-288";
            when -289 => reg3_string <= "-289";
            when -290 => reg3_string <= "-290";
            when -291 => reg3_string <= "-291";
            when -292 => reg3_string <= "-292";
            when -293 => reg3_string <= "-293";
            when -294 => reg3_string <= "-294";
            when -295 => reg3_string <= "-295";
            when -296 => reg3_string <= "-296";
            when -297 => reg3_string <= "-297";
            when -298 => reg3_string <= "-298";
            when -299 => reg3_string <= "-299";
            when -300 => reg3_string <= "-300";
            when -301 => reg3_string <= "-301";
            when -302 => reg3_string <= "-302";
            when -303 => reg3_string <= "-303";
            when -304 => reg3_string <= "-304";
            when -305 => reg3_string <= "-305";
            when -306 => reg3_string <= "-306";
            when -307 => reg3_string <= "-307";
            when -308 => reg3_string <= "-308";
            when -309 => reg3_string <= "-309";
            when -310 => reg3_string <= "-310";
            when -311 => reg3_string <= "-311";
            when -312 => reg3_string <= "-312";
            when -313 => reg3_string <= "-313";
            when -314 => reg3_string <= "-314";
            when -315 => reg3_string <= "-315";
            when -316 => reg3_string <= "-316";
            when -317 => reg3_string <= "-317";
            when -318 => reg3_string <= "-318";
            when -319 => reg3_string <= "-319";
            when -320 => reg3_string <= "-320";
            when -321 => reg3_string <= "-321";
            when -322 => reg3_string <= "-322";
            when -323 => reg3_string <= "-323";
            when -324 => reg3_string <= "-324";
            when -325 => reg3_string <= "-325";
            when -326 => reg3_string <= "-326";
            when -327 => reg3_string <= "-327";
            when -328 => reg3_string <= "-328";
            when -329 => reg3_string <= "-329";
            when -330 => reg3_string <= "-330";
            when -331 => reg3_string <= "-331";
            when -332 => reg3_string <= "-332";
            when -333 => reg3_string <= "-333";
            when -334 => reg3_string <= "-334";
            when -335 => reg3_string <= "-335";
            when -336 => reg3_string <= "-336";
            when -337 => reg3_string <= "-337";
            when -338 => reg3_string <= "-338";
            when -339 => reg3_string <= "-339";
            when -340 => reg3_string <= "-340";
            when -341 => reg3_string <= "-341";
            when -342 => reg3_string <= "-342";
            when -343 => reg3_string <= "-343";
            when -344 => reg3_string <= "-344";
            when -345 => reg3_string <= "-345";
            when -346 => reg3_string <= "-346";
            when -347 => reg3_string <= "-347";
            when -348 => reg3_string <= "-348";
            when -349 => reg3_string <= "-349";
            when -350 => reg3_string <= "-350";
            when -351 => reg3_string <= "-351";
            when -352 => reg3_string <= "-352";
            when -353 => reg3_string <= "-353";
            when -354 => reg3_string <= "-354";
            when -355 => reg3_string <= "-355";
            when -356 => reg3_string <= "-356";
            when -357 => reg3_string <= "-357";
            when -358 => reg3_string <= "-358";
            when -359 => reg3_string <= "-359";
            when -360 => reg3_string <= "-360";
            when -361 => reg3_string <= "-361";
            when -362 => reg3_string <= "-362";
            when -363 => reg3_string <= "-363";
            when -364 => reg3_string <= "-364";
            when -365 => reg3_string <= "-365";
            when -366 => reg3_string <= "-366";
            when -367 => reg3_string <= "-367";
            when -368 => reg3_string <= "-368";
            when -369 => reg3_string <= "-369";
            when -370 => reg3_string <= "-370";
            when -371 => reg3_string <= "-371";
            when -372 => reg3_string <= "-372";
            when -373 => reg3_string <= "-373";
            when -374 => reg3_string <= "-374";
            when -375 => reg3_string <= "-375";
            when -376 => reg3_string <= "-376";
            when -377 => reg3_string <= "-377";
            when -378 => reg3_string <= "-378";
            when -379 => reg3_string <= "-379";
            when -380 => reg3_string <= "-380";
            when -381 => reg3_string <= "-381";
            when -382 => reg3_string <= "-382";
            when -383 => reg3_string <= "-383";
            when -384 => reg3_string <= "-384";
            when -385 => reg3_string <= "-385";
            when -386 => reg3_string <= "-386";
            when -387 => reg3_string <= "-387";
            when -388 => reg3_string <= "-388";
            when -389 => reg3_string <= "-389";
            when -390 => reg3_string <= "-390";
            when -391 => reg3_string <= "-391";
            when -392 => reg3_string <= "-392";
            when -393 => reg3_string <= "-393";
            when -394 => reg3_string <= "-394";
            when -395 => reg3_string <= "-395";
            when -396 => reg3_string <= "-396";
            when -397 => reg3_string <= "-397";
            when -398 => reg3_string <= "-398";
            when -399 => reg3_string <= "-399";
            when -400 => reg3_string <= "-400";
            when -401 => reg3_string <= "-401";
            when -402 => reg3_string <= "-402";
            when -403 => reg3_string <= "-403";
            when -404 => reg3_string <= "-404";
            when -405 => reg3_string <= "-405";
            when -406 => reg3_string <= "-406";
            when -407 => reg3_string <= "-407";
            when -408 => reg3_string <= "-408";
            when -409 => reg3_string <= "-409";
            when -410 => reg3_string <= "-410";
            when -411 => reg3_string <= "-411";
            when -412 => reg3_string <= "-412";
            when -413 => reg3_string <= "-413";
            when -414 => reg3_string <= "-414";
            when -415 => reg3_string <= "-415";
            when -416 => reg3_string <= "-416";
            when -417 => reg3_string <= "-417";
            when -418 => reg3_string <= "-418";
            when -419 => reg3_string <= "-419";
            when -420 => reg3_string <= "-420";
            when -421 => reg3_string <= "-421";
            when -422 => reg3_string <= "-422";
            when -423 => reg3_string <= "-423";
            when -424 => reg3_string <= "-424";
            when -425 => reg3_string <= "-425";
            when -426 => reg3_string <= "-426";
            when -427 => reg3_string <= "-427";
            when -428 => reg3_string <= "-428";
            when -429 => reg3_string <= "-429";
            when -430 => reg3_string <= "-430";
            when -431 => reg3_string <= "-431";
            when -432 => reg3_string <= "-432";
            when -433 => reg3_string <= "-433";
            when -434 => reg3_string <= "-434";
            when -435 => reg3_string <= "-435";
            when -436 => reg3_string <= "-436";
            when -437 => reg3_string <= "-437";
            when -438 => reg3_string <= "-438";
            when -439 => reg3_string <= "-439";
            when -440 => reg3_string <= "-440";
            when -441 => reg3_string <= "-441";
            when -442 => reg3_string <= "-442";
            when -443 => reg3_string <= "-443";
            when -444 => reg3_string <= "-444";
            when -445 => reg3_string <= "-445";
            when -446 => reg3_string <= "-446";
            when -447 => reg3_string <= "-447";
            when -448 => reg3_string <= "-448";
            when -449 => reg3_string <= "-449";
            when -450 => reg3_string <= "-450";
            when -451 => reg3_string <= "-451";
            when -452 => reg3_string <= "-452";
            when -453 => reg3_string <= "-453";
            when -454 => reg3_string <= "-454";
            when -455 => reg3_string <= "-455";
            when -456 => reg3_string <= "-456";
            when -457 => reg3_string <= "-457";
            when -458 => reg3_string <= "-458";
            when -459 => reg3_string <= "-459";
            when -460 => reg3_string <= "-460";
            when -461 => reg3_string <= "-461";
            when -462 => reg3_string <= "-462";
            when -463 => reg3_string <= "-463";
            when -464 => reg3_string <= "-464";
            when -465 => reg3_string <= "-465";
            when -466 => reg3_string <= "-466";
            when -467 => reg3_string <= "-467";
            when -468 => reg3_string <= "-468";
            when -469 => reg3_string <= "-469";
            when -470 => reg3_string <= "-470";
            when -471 => reg3_string <= "-471";
            when -472 => reg3_string <= "-472";
            when -473 => reg3_string <= "-473";
            when -474 => reg3_string <= "-474";
            when -475 => reg3_string <= "-475";
            when -476 => reg3_string <= "-476";
            when -477 => reg3_string <= "-477";
            when -478 => reg3_string <= "-478";
            when -479 => reg3_string <= "-479";
            when -480 => reg3_string <= "-480";
            when -481 => reg3_string <= "-481";
            when -482 => reg3_string <= "-482";
            when -483 => reg3_string <= "-483";
            when -484 => reg3_string <= "-484";
            when -485 => reg3_string <= "-485";
            when -486 => reg3_string <= "-486";
            when -487 => reg3_string <= "-487";
            when -488 => reg3_string <= "-488";
            when -489 => reg3_string <= "-489";
            when -490 => reg3_string <= "-490";
            when -491 => reg3_string <= "-491";
            when -492 => reg3_string <= "-492";
            when -493 => reg3_string <= "-493";
            when -494 => reg3_string <= "-494";
            when -495 => reg3_string <= "-495";
            when -496 => reg3_string <= "-496";
            when -497 => reg3_string <= "-497";
            when -498 => reg3_string <= "-498";
            when -499 => reg3_string <= "-499";
            when -500 => reg3_string <= "-500";
            when -501 => reg3_string <= "-501";
            when -502 => reg3_string <= "-502";
            when -503 => reg3_string <= "-503";
            when -504 => reg3_string <= "-504";
            when -505 => reg3_string <= "-505";
            when -506 => reg3_string <= "-506";
            when -507 => reg3_string <= "-507";
            when -508 => reg3_string <= "-508";
            when -509 => reg3_string <= "-509";
            when -510 => reg3_string <= "-510";
            when -511 => reg3_string <= "-511";
            when -512 => reg3_string <= "-512";
            when -513 => reg3_string <= "-513";
            when -514 => reg3_string <= "-514";
            when -515 => reg3_string <= "-515";
            when -516 => reg3_string <= "-516";
            when -517 => reg3_string <= "-517";
            when -518 => reg3_string <= "-518";
            when -519 => reg3_string <= "-519";
            when -520 => reg3_string <= "-520";
            when -521 => reg3_string <= "-521";
            when -522 => reg3_string <= "-522";
            when -523 => reg3_string <= "-523";
            when -524 => reg3_string <= "-524";
            when -525 => reg3_string <= "-525";
            when -526 => reg3_string <= "-526";
            when -527 => reg3_string <= "-527";
            when -528 => reg3_string <= "-528";
            when -529 => reg3_string <= "-529";
            when -530 => reg3_string <= "-530";
            when -531 => reg3_string <= "-531";
            when -532 => reg3_string <= "-532";
            when -533 => reg3_string <= "-533";
            when -534 => reg3_string <= "-534";
            when -535 => reg3_string <= "-535";
            when -536 => reg3_string <= "-536";
            when -537 => reg3_string <= "-537";
            when -538 => reg3_string <= "-538";
            when -539 => reg3_string <= "-539";
            when -540 => reg3_string <= "-540";
            when -541 => reg3_string <= "-541";
            when -542 => reg3_string <= "-542";
            when -543 => reg3_string <= "-543";
            when -544 => reg3_string <= "-544";
            when -545 => reg3_string <= "-545";
            when -546 => reg3_string <= "-546";
            when -547 => reg3_string <= "-547";
            when -548 => reg3_string <= "-548";
            when -549 => reg3_string <= "-549";
            when -550 => reg3_string <= "-550";
            when -551 => reg3_string <= "-551";
            when -552 => reg3_string <= "-552";
            when -553 => reg3_string <= "-553";
            when -554 => reg3_string <= "-554";
            when -555 => reg3_string <= "-555";
            when -556 => reg3_string <= "-556";
            when -557 => reg3_string <= "-557";
            when -558 => reg3_string <= "-558";
            when -559 => reg3_string <= "-559";
            when -560 => reg3_string <= "-560";
            when -561 => reg3_string <= "-561";
            when -562 => reg3_string <= "-562";
            when -563 => reg3_string <= "-563";
            when -564 => reg3_string <= "-564";
            when -565 => reg3_string <= "-565";
            when -566 => reg3_string <= "-566";
            when -567 => reg3_string <= "-567";
            when -568 => reg3_string <= "-568";
            when -569 => reg3_string <= "-569";
            when -570 => reg3_string <= "-570";
            when -571 => reg3_string <= "-571";
            when -572 => reg3_string <= "-572";
            when -573 => reg3_string <= "-573";
            when -574 => reg3_string <= "-574";
            when -575 => reg3_string <= "-575";
            when -576 => reg3_string <= "-576";
            when -577 => reg3_string <= "-577";
            when -578 => reg3_string <= "-578";
            when -579 => reg3_string <= "-579";
            when -580 => reg3_string <= "-580";
            when -581 => reg3_string <= "-581";
            when -582 => reg3_string <= "-582";
            when -583 => reg3_string <= "-583";
            when -584 => reg3_string <= "-584";
            when -585 => reg3_string <= "-585";
            when -586 => reg3_string <= "-586";
            when -587 => reg3_string <= "-587";
            when -588 => reg3_string <= "-588";
            when -589 => reg3_string <= "-589";
            when -590 => reg3_string <= "-590";
            when -591 => reg3_string <= "-591";
            when -592 => reg3_string <= "-592";
            when -593 => reg3_string <= "-593";
            when -594 => reg3_string <= "-594";
            when -595 => reg3_string <= "-595";
            when -596 => reg3_string <= "-596";
            when -597 => reg3_string <= "-597";
            when -598 => reg3_string <= "-598";
            when -599 => reg3_string <= "-599";
            when -600 => reg3_string <= "-600";
            when -601 => reg3_string <= "-601";
            when -602 => reg3_string <= "-602";
            when -603 => reg3_string <= "-603";
            when -604 => reg3_string <= "-604";
            when -605 => reg3_string <= "-605";
            when -606 => reg3_string <= "-606";
            when -607 => reg3_string <= "-607";
            when -608 => reg3_string <= "-608";
            when -609 => reg3_string <= "-609";
            when -610 => reg3_string <= "-610";
            when -611 => reg3_string <= "-611";
            when -612 => reg3_string <= "-612";
            when -613 => reg3_string <= "-613";
            when -614 => reg3_string <= "-614";
            when -615 => reg3_string <= "-615";
            when -616 => reg3_string <= "-616";
            when -617 => reg3_string <= "-617";
            when -618 => reg3_string <= "-618";
            when -619 => reg3_string <= "-619";
            when -620 => reg3_string <= "-620";
            when -621 => reg3_string <= "-621";
            when -622 => reg3_string <= "-622";
            when -623 => reg3_string <= "-623";
            when -624 => reg3_string <= "-624";
            when -625 => reg3_string <= "-625";
            when -626 => reg3_string <= "-626";
            when -627 => reg3_string <= "-627";
            when -628 => reg3_string <= "-628";
            when -629 => reg3_string <= "-629";
            when -630 => reg3_string <= "-630";
            when -631 => reg3_string <= "-631";
            when -632 => reg3_string <= "-632";
            when -633 => reg3_string <= "-633";
            when -634 => reg3_string <= "-634";
            when -635 => reg3_string <= "-635";
            when -636 => reg3_string <= "-636";
            when -637 => reg3_string <= "-637";
            when -638 => reg3_string <= "-638";
            when -639 => reg3_string <= "-639";
            when -640 => reg3_string <= "-640";
            when -641 => reg3_string <= "-641";
            when -642 => reg3_string <= "-642";
            when -643 => reg3_string <= "-643";
            when -644 => reg3_string <= "-644";
            when -645 => reg3_string <= "-645";
            when -646 => reg3_string <= "-646";
            when -647 => reg3_string <= "-647";
            when -648 => reg3_string <= "-648";
            when -649 => reg3_string <= "-649";
            when -650 => reg3_string <= "-650";
            when -651 => reg3_string <= "-651";
            when -652 => reg3_string <= "-652";
            when -653 => reg3_string <= "-653";
            when -654 => reg3_string <= "-654";
            when -655 => reg3_string <= "-655";
            when -656 => reg3_string <= "-656";
            when -657 => reg3_string <= "-657";
            when -658 => reg3_string <= "-658";
            when -659 => reg3_string <= "-659";
            when -660 => reg3_string <= "-660";
            when -661 => reg3_string <= "-661";
            when -662 => reg3_string <= "-662";
            when -663 => reg3_string <= "-663";
            when -664 => reg3_string <= "-664";
            when -665 => reg3_string <= "-665";
            when -666 => reg3_string <= "-666";
            when -667 => reg3_string <= "-667";
            when -668 => reg3_string <= "-668";
            when -669 => reg3_string <= "-669";
            when -670 => reg3_string <= "-670";
            when -671 => reg3_string <= "-671";
            when -672 => reg3_string <= "-672";
            when -673 => reg3_string <= "-673";
            when -674 => reg3_string <= "-674";
            when -675 => reg3_string <= "-675";
            when -676 => reg3_string <= "-676";
            when -677 => reg3_string <= "-677";
            when -678 => reg3_string <= "-678";
            when -679 => reg3_string <= "-679";
            when -680 => reg3_string <= "-680";
            when -681 => reg3_string <= "-681";
            when -682 => reg3_string <= "-682";
            when -683 => reg3_string <= "-683";
            when -684 => reg3_string <= "-684";
            when -685 => reg3_string <= "-685";
            when -686 => reg3_string <= "-686";
            when -687 => reg3_string <= "-687";
            when -688 => reg3_string <= "-688";
            when -689 => reg3_string <= "-689";
            when -690 => reg3_string <= "-690";
            when -691 => reg3_string <= "-691";
            when -692 => reg3_string <= "-692";
            when -693 => reg3_string <= "-693";
            when -694 => reg3_string <= "-694";
            when -695 => reg3_string <= "-695";
            when -696 => reg3_string <= "-696";
            when -697 => reg3_string <= "-697";
            when -698 => reg3_string <= "-698";
            when -699 => reg3_string <= "-699";
            when -700 => reg3_string <= "-700";
            when -701 => reg3_string <= "-701";
            when -702 => reg3_string <= "-702";
            when -703 => reg3_string <= "-703";
            when -704 => reg3_string <= "-704";
            when -705 => reg3_string <= "-705";
            when -706 => reg3_string <= "-706";
            when -707 => reg3_string <= "-707";
            when -708 => reg3_string <= "-708";
            when -709 => reg3_string <= "-709";
            when -710 => reg3_string <= "-710";
            when -711 => reg3_string <= "-711";
            when -712 => reg3_string <= "-712";
            when -713 => reg3_string <= "-713";
            when -714 => reg3_string <= "-714";
            when -715 => reg3_string <= "-715";
            when -716 => reg3_string <= "-716";
            when -717 => reg3_string <= "-717";
            when -718 => reg3_string <= "-718";
            when -719 => reg3_string <= "-719";
            when -720 => reg3_string <= "-720";
            when -721 => reg3_string <= "-721";
            when -722 => reg3_string <= "-722";
            when -723 => reg3_string <= "-723";
            when -724 => reg3_string <= "-724";
            when -725 => reg3_string <= "-725";
            when -726 => reg3_string <= "-726";
            when -727 => reg3_string <= "-727";
            when -728 => reg3_string <= "-728";
            when -729 => reg3_string <= "-729";
            when -730 => reg3_string <= "-730";
            when -731 => reg3_string <= "-731";
            when -732 => reg3_string <= "-732";
            when -733 => reg3_string <= "-733";
            when -734 => reg3_string <= "-734";
            when -735 => reg3_string <= "-735";
            when -736 => reg3_string <= "-736";
            when -737 => reg3_string <= "-737";
            when -738 => reg3_string <= "-738";
            when -739 => reg3_string <= "-739";
            when -740 => reg3_string <= "-740";
            when -741 => reg3_string <= "-741";
            when -742 => reg3_string <= "-742";
            when -743 => reg3_string <= "-743";
            when -744 => reg3_string <= "-744";
            when -745 => reg3_string <= "-745";
            when -746 => reg3_string <= "-746";
            when -747 => reg3_string <= "-747";
            when -748 => reg3_string <= "-748";
            when -749 => reg3_string <= "-749";
            when -750 => reg3_string <= "-750";
            when -751 => reg3_string <= "-751";
            when -752 => reg3_string <= "-752";
            when -753 => reg3_string <= "-753";
            when -754 => reg3_string <= "-754";
            when -755 => reg3_string <= "-755";
            when -756 => reg3_string <= "-756";
            when -757 => reg3_string <= "-757";
            when -758 => reg3_string <= "-758";
            when -759 => reg3_string <= "-759";
            when -760 => reg3_string <= "-760";
            when -761 => reg3_string <= "-761";
            when -762 => reg3_string <= "-762";
            when -763 => reg3_string <= "-763";
            when -764 => reg3_string <= "-764";
            when -765 => reg3_string <= "-765";
            when -766 => reg3_string <= "-766";
            when -767 => reg3_string <= "-767";
            when -768 => reg3_string <= "-768";
            when -769 => reg3_string <= "-769";
            when -770 => reg3_string <= "-770";
            when -771 => reg3_string <= "-771";
            when -772 => reg3_string <= "-772";
            when -773 => reg3_string <= "-773";
            when -774 => reg3_string <= "-774";
            when -775 => reg3_string <= "-775";
            when -776 => reg3_string <= "-776";
            when -777 => reg3_string <= "-777";
            when -778 => reg3_string <= "-778";
            when -779 => reg3_string <= "-779";
            when -780 => reg3_string <= "-780";
            when -781 => reg3_string <= "-781";
            when -782 => reg3_string <= "-782";
            when -783 => reg3_string <= "-783";
            when -784 => reg3_string <= "-784";
            when -785 => reg3_string <= "-785";
            when -786 => reg3_string <= "-786";
            when -787 => reg3_string <= "-787";
            when -788 => reg3_string <= "-788";
            when -789 => reg3_string <= "-789";
            when -790 => reg3_string <= "-790";
            when -791 => reg3_string <= "-791";
            when -792 => reg3_string <= "-792";
            when -793 => reg3_string <= "-793";
            when -794 => reg3_string <= "-794";
            when -795 => reg3_string <= "-795";
            when -796 => reg3_string <= "-796";
            when -797 => reg3_string <= "-797";
            when -798 => reg3_string <= "-798";
            when -799 => reg3_string <= "-799";
            when -800 => reg3_string <= "-800";
            when -801 => reg3_string <= "-801";
            when -802 => reg3_string <= "-802";
            when -803 => reg3_string <= "-803";
            when -804 => reg3_string <= "-804";
            when -805 => reg3_string <= "-805";
            when -806 => reg3_string <= "-806";
            when -807 => reg3_string <= "-807";
            when -808 => reg3_string <= "-808";
            when -809 => reg3_string <= "-809";
            when -810 => reg3_string <= "-810";
            when -811 => reg3_string <= "-811";
            when -812 => reg3_string <= "-812";
            when -813 => reg3_string <= "-813";
            when -814 => reg3_string <= "-814";
            when -815 => reg3_string <= "-815";
            when -816 => reg3_string <= "-816";
            when -817 => reg3_string <= "-817";
            when -818 => reg3_string <= "-818";
            when -819 => reg3_string <= "-819";
            when -820 => reg3_string <= "-820";
            when -821 => reg3_string <= "-821";
            when -822 => reg3_string <= "-822";
            when -823 => reg3_string <= "-823";
            when -824 => reg3_string <= "-824";
            when -825 => reg3_string <= "-825";
            when -826 => reg3_string <= "-826";
            when -827 => reg3_string <= "-827";
            when -828 => reg3_string <= "-828";
            when -829 => reg3_string <= "-829";
            when -830 => reg3_string <= "-830";
            when -831 => reg3_string <= "-831";
            when -832 => reg3_string <= "-832";
            when -833 => reg3_string <= "-833";
            when -834 => reg3_string <= "-834";
            when -835 => reg3_string <= "-835";
            when -836 => reg3_string <= "-836";
            when -837 => reg3_string <= "-837";
            when -838 => reg3_string <= "-838";
            when -839 => reg3_string <= "-839";
            when -840 => reg3_string <= "-840";
            when -841 => reg3_string <= "-841";
            when -842 => reg3_string <= "-842";
            when -843 => reg3_string <= "-843";
            when -844 => reg3_string <= "-844";
            when -845 => reg3_string <= "-845";
            when -846 => reg3_string <= "-846";
            when -847 => reg3_string <= "-847";
            when -848 => reg3_string <= "-848";
            when -849 => reg3_string <= "-849";
            when -850 => reg3_string <= "-850";
            when -851 => reg3_string <= "-851";
            when -852 => reg3_string <= "-852";
            when -853 => reg3_string <= "-853";
            when -854 => reg3_string <= "-854";
            when -855 => reg3_string <= "-855";
            when -856 => reg3_string <= "-856";
            when -857 => reg3_string <= "-857";
            when -858 => reg3_string <= "-858";
            when -859 => reg3_string <= "-859";
            when -860 => reg3_string <= "-860";
            when -861 => reg3_string <= "-861";
            when -862 => reg3_string <= "-862";
            when -863 => reg3_string <= "-863";
            when -864 => reg3_string <= "-864";
            when -865 => reg3_string <= "-865";
            when -866 => reg3_string <= "-866";
            when -867 => reg3_string <= "-867";
            when -868 => reg3_string <= "-868";
            when -869 => reg3_string <= "-869";
            when -870 => reg3_string <= "-870";
            when -871 => reg3_string <= "-871";
            when -872 => reg3_string <= "-872";
            when -873 => reg3_string <= "-873";
            when -874 => reg3_string <= "-874";
            when -875 => reg3_string <= "-875";
            when -876 => reg3_string <= "-876";
            when -877 => reg3_string <= "-877";
            when -878 => reg3_string <= "-878";
            when -879 => reg3_string <= "-879";
            when -880 => reg3_string <= "-880";
            when -881 => reg3_string <= "-881";
            when -882 => reg3_string <= "-882";
            when -883 => reg3_string <= "-883";
            when -884 => reg3_string <= "-884";
            when -885 => reg3_string <= "-885";
            when -886 => reg3_string <= "-886";
            when -887 => reg3_string <= "-887";
            when -888 => reg3_string <= "-888";
            when -889 => reg3_string <= "-889";
            when -890 => reg3_string <= "-890";
            when -891 => reg3_string <= "-891";
            when -892 => reg3_string <= "-892";
            when -893 => reg3_string <= "-893";
            when -894 => reg3_string <= "-894";
            when -895 => reg3_string <= "-895";
            when -896 => reg3_string <= "-896";
            when -897 => reg3_string <= "-897";
            when -898 => reg3_string <= "-898";
            when -899 => reg3_string <= "-899";
            when -900 => reg3_string <= "-900";
            when -901 => reg3_string <= "-901";
            when -902 => reg3_string <= "-902";
            when -903 => reg3_string <= "-903";
            when -904 => reg3_string <= "-904";
            when -905 => reg3_string <= "-905";
            when -906 => reg3_string <= "-906";
            when -907 => reg3_string <= "-907";
            when -908 => reg3_string <= "-908";
            when -909 => reg3_string <= "-909";
            when -910 => reg3_string <= "-910";
            when -911 => reg3_string <= "-911";
            when -912 => reg3_string <= "-912";
            when -913 => reg3_string <= "-913";
            when -914 => reg3_string <= "-914";
            when -915 => reg3_string <= "-915";
            when -916 => reg3_string <= "-916";
            when -917 => reg3_string <= "-917";
            when -918 => reg3_string <= "-918";
            when -919 => reg3_string <= "-919";
            when -920 => reg3_string <= "-920";
            when -921 => reg3_string <= "-921";
            when -922 => reg3_string <= "-922";
            when -923 => reg3_string <= "-923";
            when -924 => reg3_string <= "-924";
            when -925 => reg3_string <= "-925";
            when -926 => reg3_string <= "-926";
            when -927 => reg3_string <= "-927";
            when -928 => reg3_string <= "-928";
            when -929 => reg3_string <= "-929";
            when -930 => reg3_string <= "-930";
            when -931 => reg3_string <= "-931";
            when -932 => reg3_string <= "-932";
            when -933 => reg3_string <= "-933";
            when -934 => reg3_string <= "-934";
            when -935 => reg3_string <= "-935";
            when -936 => reg3_string <= "-936";
            when -937 => reg3_string <= "-937";
            when -938 => reg3_string <= "-938";
            when -939 => reg3_string <= "-939";
            when -940 => reg3_string <= "-940";
            when -941 => reg3_string <= "-941";
            when -942 => reg3_string <= "-942";
            when -943 => reg3_string <= "-943";
            when -944 => reg3_string <= "-944";
            when -945 => reg3_string <= "-945";
            when -946 => reg3_string <= "-946";
            when -947 => reg3_string <= "-947";
            when -948 => reg3_string <= "-948";
            when -949 => reg3_string <= "-949";
            when -950 => reg3_string <= "-950";
            when -951 => reg3_string <= "-951";
            when -952 => reg3_string <= "-952";
            when -953 => reg3_string <= "-953";
            when -954 => reg3_string <= "-954";
            when -955 => reg3_string <= "-955";
            when -956 => reg3_string <= "-956";
            when -957 => reg3_string <= "-957";
            when -958 => reg3_string <= "-958";
            when -959 => reg3_string <= "-959";
            when -960 => reg3_string <= "-960";
            when -961 => reg3_string <= "-961";
            when -962 => reg3_string <= "-962";
            when -963 => reg3_string <= "-963";
            when -964 => reg3_string <= "-964";
            when -965 => reg3_string <= "-965";
            when -966 => reg3_string <= "-966";
            when -967 => reg3_string <= "-967";
            when -968 => reg3_string <= "-968";
            when -969 => reg3_string <= "-969";
            when -970 => reg3_string <= "-970";
            when -971 => reg3_string <= "-971";
            when -972 => reg3_string <= "-972";
            when -973 => reg3_string <= "-973";
            when -974 => reg3_string <= "-974";
            when -975 => reg3_string <= "-975";
            when -976 => reg3_string <= "-976";
            when -977 => reg3_string <= "-977";
            when -978 => reg3_string <= "-978";
            when -979 => reg3_string <= "-979";
            when -980 => reg3_string <= "-980";
            when -981 => reg3_string <= "-981";
            when -982 => reg3_string <= "-982";
            when -983 => reg3_string <= "-983";
            when -984 => reg3_string <= "-984";
            when -985 => reg3_string <= "-985";
            when -986 => reg3_string <= "-986";
            when -987 => reg3_string <= "-987";
            when -988 => reg3_string <= "-988";
            when -989 => reg3_string <= "-989";
            when -990 => reg3_string <= "-990";
            when -991 => reg3_string <= "-991";
            when -992 => reg3_string <= "-992";
            when -993 => reg3_string <= "-993";
            when -994 => reg3_string <= "-994";
            when -995 => reg3_string <= "-995";
            when -996 => reg3_string <= "-996";
            when -997 => reg3_string <= "-997";
            when -998 => reg3_string <= "-998";
            when -999 => reg3_string <= "-999";
            when others => reg3_string <= "    ";
        end case;
        
        case (reg2_int) is 
        when 999 => reg2_string <= " 999";
        when 998 => reg2_string <= " 998";
        when 997 => reg2_string <= " 997";
        when 996 => reg2_string <= " 996";
        when 995 => reg2_string <= " 995";
        when 994 => reg2_string <= " 994";
        when 993 => reg2_string <= " 993";
        when 992 => reg2_string <= " 992";
        when 991 => reg2_string <= " 991";
        when 990 => reg2_string <= " 990";
        when 989 => reg2_string <= " 989";
        when 988 => reg2_string <= " 988";
        when 987 => reg2_string <= " 987";
        when 986 => reg2_string <= " 986";
        when 985 => reg2_string <= " 985";
        when 984 => reg2_string <= " 984";
        when 983 => reg2_string <= " 983";
        when 982 => reg2_string <= " 982";
        when 981 => reg2_string <= " 981";
        when 980 => reg2_string <= " 980";
        when 979 => reg2_string <= " 979";
        when 978 => reg2_string <= " 978";
        when 977 => reg2_string <= " 977";
        when 976 => reg2_string <= " 976";
        when 975 => reg2_string <= " 975";
        when 974 => reg2_string <= " 974";
        when 973 => reg2_string <= " 973";
        when 972 => reg2_string <= " 972";
        when 971 => reg2_string <= " 971";
        when 970 => reg2_string <= " 970";
        when 969 => reg2_string <= " 969";
        when 968 => reg2_string <= " 968";
        when 967 => reg2_string <= " 967";
        when 966 => reg2_string <= " 966";
        when 965 => reg2_string <= " 965";
        when 964 => reg2_string <= " 964";
        when 963 => reg2_string <= " 963";
        when 962 => reg2_string <= " 962";
        when 961 => reg2_string <= " 961";
        when 960 => reg2_string <= " 960";
        when 959 => reg2_string <= " 959";
        when 958 => reg2_string <= " 958";
        when 957 => reg2_string <= " 957";
        when 956 => reg2_string <= " 956";
        when 955 => reg2_string <= " 955";
        when 954 => reg2_string <= " 954";
        when 953 => reg2_string <= " 953";
        when 952 => reg2_string <= " 952";
        when 951 => reg2_string <= " 951";
        when 950 => reg2_string <= " 950";
        when 949 => reg2_string <= " 949";
        when 948 => reg2_string <= " 948";
        when 947 => reg2_string <= " 947";
        when 946 => reg2_string <= " 946";
        when 945 => reg2_string <= " 945";
        when 944 => reg2_string <= " 944";
        when 943 => reg2_string <= " 943";
        when 942 => reg2_string <= " 942";
        when 941 => reg2_string <= " 941";
        when 940 => reg2_string <= " 940";
        when 939 => reg2_string <= " 939";
        when 938 => reg2_string <= " 938";
        when 937 => reg2_string <= " 937";
        when 936 => reg2_string <= " 936";
        when 935 => reg2_string <= " 935";
        when 934 => reg2_string <= " 934";
        when 933 => reg2_string <= " 933";
        when 932 => reg2_string <= " 932";
        when 931 => reg2_string <= " 931";
        when 930 => reg2_string <= " 930";
        when 929 => reg2_string <= " 929";
        when 928 => reg2_string <= " 928";
        when 927 => reg2_string <= " 927";
        when 926 => reg2_string <= " 926";
        when 925 => reg2_string <= " 925";
        when 924 => reg2_string <= " 924";
        when 923 => reg2_string <= " 923";
        when 922 => reg2_string <= " 922";
        when 921 => reg2_string <= " 921";
        when 920 => reg2_string <= " 920";
        when 919 => reg2_string <= " 919";
        when 918 => reg2_string <= " 918";
        when 917 => reg2_string <= " 917";
        when 916 => reg2_string <= " 916";
        when 915 => reg2_string <= " 915";
        when 914 => reg2_string <= " 914";
        when 913 => reg2_string <= " 913";
        when 912 => reg2_string <= " 912";
        when 911 => reg2_string <= " 911";
        when 910 => reg2_string <= " 910";
        when 909 => reg2_string <= " 909";
        when 908 => reg2_string <= " 908";
        when 907 => reg2_string <= " 907";
        when 906 => reg2_string <= " 906";
        when 905 => reg2_string <= " 905";
        when 904 => reg2_string <= " 904";
        when 903 => reg2_string <= " 903";
        when 902 => reg2_string <= " 902";
        when 901 => reg2_string <= " 901";
        when 900 => reg2_string <= " 900";
        when 899 => reg2_string <= " 899";
        when 898 => reg2_string <= " 898";
        when 897 => reg2_string <= " 897";
        when 896 => reg2_string <= " 896";
        when 895 => reg2_string <= " 895";
        when 894 => reg2_string <= " 894";
        when 893 => reg2_string <= " 893";
        when 892 => reg2_string <= " 892";
        when 891 => reg2_string <= " 891";
        when 890 => reg2_string <= " 890";
        when 889 => reg2_string <= " 889";
        when 888 => reg2_string <= " 888";
        when 887 => reg2_string <= " 887";
        when 886 => reg2_string <= " 886";
        when 885 => reg2_string <= " 885";
        when 884 => reg2_string <= " 884";
        when 883 => reg2_string <= " 883";
        when 882 => reg2_string <= " 882";
        when 881 => reg2_string <= " 881";
        when 880 => reg2_string <= " 880";
        when 879 => reg2_string <= " 879";
        when 878 => reg2_string <= " 878";
        when 877 => reg2_string <= " 877";
        when 876 => reg2_string <= " 876";
        when 875 => reg2_string <= " 875";
        when 874 => reg2_string <= " 874";
        when 873 => reg2_string <= " 873";
        when 872 => reg2_string <= " 872";
        when 871 => reg2_string <= " 871";
        when 870 => reg2_string <= " 870";
        when 869 => reg2_string <= " 869";
        when 868 => reg2_string <= " 868";
        when 867 => reg2_string <= " 867";
        when 866 => reg2_string <= " 866";
        when 865 => reg2_string <= " 865";
        when 864 => reg2_string <= " 864";
        when 863 => reg2_string <= " 863";
        when 862 => reg2_string <= " 862";
        when 861 => reg2_string <= " 861";
        when 860 => reg2_string <= " 860";
        when 859 => reg2_string <= " 859";
        when 858 => reg2_string <= " 858";
        when 857 => reg2_string <= " 857";
        when 856 => reg2_string <= " 856";
        when 855 => reg2_string <= " 855";
        when 854 => reg2_string <= " 854";
        when 853 => reg2_string <= " 853";
        when 852 => reg2_string <= " 852";
        when 851 => reg2_string <= " 851";
        when 850 => reg2_string <= " 850";
        when 849 => reg2_string <= " 849";
        when 848 => reg2_string <= " 848";
        when 847 => reg2_string <= " 847";
        when 846 => reg2_string <= " 846";
        when 845 => reg2_string <= " 845";
        when 844 => reg2_string <= " 844";
        when 843 => reg2_string <= " 843";
        when 842 => reg2_string <= " 842";
        when 841 => reg2_string <= " 841";
        when 840 => reg2_string <= " 840";
        when 839 => reg2_string <= " 839";
        when 838 => reg2_string <= " 838";
        when 837 => reg2_string <= " 837";
        when 836 => reg2_string <= " 836";
        when 835 => reg2_string <= " 835";
        when 834 => reg2_string <= " 834";
        when 833 => reg2_string <= " 833";
        when 832 => reg2_string <= " 832";
        when 831 => reg2_string <= " 831";
        when 830 => reg2_string <= " 830";
        when 829 => reg2_string <= " 829";
        when 828 => reg2_string <= " 828";
        when 827 => reg2_string <= " 827";
        when 826 => reg2_string <= " 826";
        when 825 => reg2_string <= " 825";
        when 824 => reg2_string <= " 824";
        when 823 => reg2_string <= " 823";
        when 822 => reg2_string <= " 822";
        when 821 => reg2_string <= " 821";
        when 820 => reg2_string <= " 820";
        when 819 => reg2_string <= " 819";
        when 818 => reg2_string <= " 818";
        when 817 => reg2_string <= " 817";
        when 816 => reg2_string <= " 816";
        when 815 => reg2_string <= " 815";
        when 814 => reg2_string <= " 814";
        when 813 => reg2_string <= " 813";
        when 812 => reg2_string <= " 812";
        when 811 => reg2_string <= " 811";
        when 810 => reg2_string <= " 810";
        when 809 => reg2_string <= " 809";
        when 808 => reg2_string <= " 808";
        when 807 => reg2_string <= " 807";
        when 806 => reg2_string <= " 806";
        when 805 => reg2_string <= " 805";
        when 804 => reg2_string <= " 804";
        when 803 => reg2_string <= " 803";
        when 802 => reg2_string <= " 802";
        when 801 => reg2_string <= " 801";
        when 800 => reg2_string <= " 800";
        when 799 => reg2_string <= " 799";
        when 798 => reg2_string <= " 798";
        when 797 => reg2_string <= " 797";
        when 796 => reg2_string <= " 796";
        when 795 => reg2_string <= " 795";
        when 794 => reg2_string <= " 794";
        when 793 => reg2_string <= " 793";
        when 792 => reg2_string <= " 792";
        when 791 => reg2_string <= " 791";
        when 790 => reg2_string <= " 790";
        when 789 => reg2_string <= " 789";
        when 788 => reg2_string <= " 788";
        when 787 => reg2_string <= " 787";
        when 786 => reg2_string <= " 786";
        when 785 => reg2_string <= " 785";
        when 784 => reg2_string <= " 784";
        when 783 => reg2_string <= " 783";
        when 782 => reg2_string <= " 782";
        when 781 => reg2_string <= " 781";
        when 780 => reg2_string <= " 780";
        when 779 => reg2_string <= " 779";
        when 778 => reg2_string <= " 778";
        when 777 => reg2_string <= " 777";
        when 776 => reg2_string <= " 776";
        when 775 => reg2_string <= " 775";
        when 774 => reg2_string <= " 774";
        when 773 => reg2_string <= " 773";
        when 772 => reg2_string <= " 772";
        when 771 => reg2_string <= " 771";
        when 770 => reg2_string <= " 770";
        when 769 => reg2_string <= " 769";
        when 768 => reg2_string <= " 768";
        when 767 => reg2_string <= " 767";
        when 766 => reg2_string <= " 766";
        when 765 => reg2_string <= " 765";
        when 764 => reg2_string <= " 764";
        when 763 => reg2_string <= " 763";
        when 762 => reg2_string <= " 762";
        when 761 => reg2_string <= " 761";
        when 760 => reg2_string <= " 760";
        when 759 => reg2_string <= " 759";
        when 758 => reg2_string <= " 758";
        when 757 => reg2_string <= " 757";
        when 756 => reg2_string <= " 756";
        when 755 => reg2_string <= " 755";
        when 754 => reg2_string <= " 754";
        when 753 => reg2_string <= " 753";
        when 752 => reg2_string <= " 752";
        when 751 => reg2_string <= " 751";
        when 750 => reg2_string <= " 750";
        when 749 => reg2_string <= " 749";
        when 748 => reg2_string <= " 748";
        when 747 => reg2_string <= " 747";
        when 746 => reg2_string <= " 746";
        when 745 => reg2_string <= " 745";
        when 744 => reg2_string <= " 744";
        when 743 => reg2_string <= " 743";
        when 742 => reg2_string <= " 742";
        when 741 => reg2_string <= " 741";
        when 740 => reg2_string <= " 740";
        when 739 => reg2_string <= " 739";
        when 738 => reg2_string <= " 738";
        when 737 => reg2_string <= " 737";
        when 736 => reg2_string <= " 736";
        when 735 => reg2_string <= " 735";
        when 734 => reg2_string <= " 734";
        when 733 => reg2_string <= " 733";
        when 732 => reg2_string <= " 732";
        when 731 => reg2_string <= " 731";
        when 730 => reg2_string <= " 730";
        when 729 => reg2_string <= " 729";
        when 728 => reg2_string <= " 728";
        when 727 => reg2_string <= " 727";
        when 726 => reg2_string <= " 726";
        when 725 => reg2_string <= " 725";
        when 724 => reg2_string <= " 724";
        when 723 => reg2_string <= " 723";
        when 722 => reg2_string <= " 722";
        when 721 => reg2_string <= " 721";
        when 720 => reg2_string <= " 720";
        when 719 => reg2_string <= " 719";
        when 718 => reg2_string <= " 718";
        when 717 => reg2_string <= " 717";
        when 716 => reg2_string <= " 716";
        when 715 => reg2_string <= " 715";
        when 714 => reg2_string <= " 714";
        when 713 => reg2_string <= " 713";
        when 712 => reg2_string <= " 712";
        when 711 => reg2_string <= " 711";
        when 710 => reg2_string <= " 710";
        when 709 => reg2_string <= " 709";
        when 708 => reg2_string <= " 708";
        when 707 => reg2_string <= " 707";
        when 706 => reg2_string <= " 706";
        when 705 => reg2_string <= " 705";
        when 704 => reg2_string <= " 704";
        when 703 => reg2_string <= " 703";
        when 702 => reg2_string <= " 702";
        when 701 => reg2_string <= " 701";
        when 700 => reg2_string <= " 700";
        when 699 => reg2_string <= " 699";
        when 698 => reg2_string <= " 698";
        when 697 => reg2_string <= " 697";
        when 696 => reg2_string <= " 696";
        when 695 => reg2_string <= " 695";
        when 694 => reg2_string <= " 694";
        when 693 => reg2_string <= " 693";
        when 692 => reg2_string <= " 692";
        when 691 => reg2_string <= " 691";
        when 690 => reg2_string <= " 690";
        when 689 => reg2_string <= " 689";
        when 688 => reg2_string <= " 688";
        when 687 => reg2_string <= " 687";
        when 686 => reg2_string <= " 686";
        when 685 => reg2_string <= " 685";
        when 684 => reg2_string <= " 684";
        when 683 => reg2_string <= " 683";
        when 682 => reg2_string <= " 682";
        when 681 => reg2_string <= " 681";
        when 680 => reg2_string <= " 680";
        when 679 => reg2_string <= " 679";
        when 678 => reg2_string <= " 678";
        when 677 => reg2_string <= " 677";
        when 676 => reg2_string <= " 676";
        when 675 => reg2_string <= " 675";
        when 674 => reg2_string <= " 674";
        when 673 => reg2_string <= " 673";
        when 672 => reg2_string <= " 672";
        when 671 => reg2_string <= " 671";
        when 670 => reg2_string <= " 670";
        when 669 => reg2_string <= " 669";
        when 668 => reg2_string <= " 668";
        when 667 => reg2_string <= " 667";
        when 666 => reg2_string <= " 666";
        when 665 => reg2_string <= " 665";
        when 664 => reg2_string <= " 664";
        when 663 => reg2_string <= " 663";
        when 662 => reg2_string <= " 662";
        when 661 => reg2_string <= " 661";
        when 660 => reg2_string <= " 660";
        when 659 => reg2_string <= " 659";
        when 658 => reg2_string <= " 658";
        when 657 => reg2_string <= " 657";
        when 656 => reg2_string <= " 656";
        when 655 => reg2_string <= " 655";
        when 654 => reg2_string <= " 654";
        when 653 => reg2_string <= " 653";
        when 652 => reg2_string <= " 652";
        when 651 => reg2_string <= " 651";
        when 650 => reg2_string <= " 650";
        when 649 => reg2_string <= " 649";
        when 648 => reg2_string <= " 648";
        when 647 => reg2_string <= " 647";
        when 646 => reg2_string <= " 646";
        when 645 => reg2_string <= " 645";
        when 644 => reg2_string <= " 644";
        when 643 => reg2_string <= " 643";
        when 642 => reg2_string <= " 642";
        when 641 => reg2_string <= " 641";
        when 640 => reg2_string <= " 640";
        when 639 => reg2_string <= " 639";
        when 638 => reg2_string <= " 638";
        when 637 => reg2_string <= " 637";
        when 636 => reg2_string <= " 636";
        when 635 => reg2_string <= " 635";
        when 634 => reg2_string <= " 634";
        when 633 => reg2_string <= " 633";
        when 632 => reg2_string <= " 632";
        when 631 => reg2_string <= " 631";
        when 630 => reg2_string <= " 630";
        when 629 => reg2_string <= " 629";
        when 628 => reg2_string <= " 628";
        when 627 => reg2_string <= " 627";
        when 626 => reg2_string <= " 626";
        when 625 => reg2_string <= " 625";
        when 624 => reg2_string <= " 624";
        when 623 => reg2_string <= " 623";
        when 622 => reg2_string <= " 622";
        when 621 => reg2_string <= " 621";
        when 620 => reg2_string <= " 620";
        when 619 => reg2_string <= " 619";
        when 618 => reg2_string <= " 618";
        when 617 => reg2_string <= " 617";
        when 616 => reg2_string <= " 616";
        when 615 => reg2_string <= " 615";
        when 614 => reg2_string <= " 614";
        when 613 => reg2_string <= " 613";
        when 612 => reg2_string <= " 612";
        when 611 => reg2_string <= " 611";
        when 610 => reg2_string <= " 610";
        when 609 => reg2_string <= " 609";
        when 608 => reg2_string <= " 608";
        when 607 => reg2_string <= " 607";
        when 606 => reg2_string <= " 606";
        when 605 => reg2_string <= " 605";
        when 604 => reg2_string <= " 604";
        when 603 => reg2_string <= " 603";
        when 602 => reg2_string <= " 602";
        when 601 => reg2_string <= " 601";
        when 600 => reg2_string <= " 600";
        when 599 => reg2_string <= " 599";
        when 598 => reg2_string <= " 598";
        when 597 => reg2_string <= " 597";
        when 596 => reg2_string <= " 596";
        when 595 => reg2_string <= " 595";
        when 594 => reg2_string <= " 594";
        when 593 => reg2_string <= " 593";
        when 592 => reg2_string <= " 592";
        when 591 => reg2_string <= " 591";
        when 590 => reg2_string <= " 590";
        when 589 => reg2_string <= " 589";
        when 588 => reg2_string <= " 588";
        when 587 => reg2_string <= " 587";
        when 586 => reg2_string <= " 586";
        when 585 => reg2_string <= " 585";
        when 584 => reg2_string <= " 584";
        when 583 => reg2_string <= " 583";
        when 582 => reg2_string <= " 582";
        when 581 => reg2_string <= " 581";
        when 580 => reg2_string <= " 580";
        when 579 => reg2_string <= " 579";
        when 578 => reg2_string <= " 578";
        when 577 => reg2_string <= " 577";
        when 576 => reg2_string <= " 576";
        when 575 => reg2_string <= " 575";
        when 574 => reg2_string <= " 574";
        when 573 => reg2_string <= " 573";
        when 572 => reg2_string <= " 572";
        when 571 => reg2_string <= " 571";
        when 570 => reg2_string <= " 570";
        when 569 => reg2_string <= " 569";
        when 568 => reg2_string <= " 568";
        when 567 => reg2_string <= " 567";
        when 566 => reg2_string <= " 566";
        when 565 => reg2_string <= " 565";
        when 564 => reg2_string <= " 564";
        when 563 => reg2_string <= " 563";
        when 562 => reg2_string <= " 562";
        when 561 => reg2_string <= " 561";
        when 560 => reg2_string <= " 560";
        when 559 => reg2_string <= " 559";
        when 558 => reg2_string <= " 558";
        when 557 => reg2_string <= " 557";
        when 556 => reg2_string <= " 556";
        when 555 => reg2_string <= " 555";
        when 554 => reg2_string <= " 554";
        when 553 => reg2_string <= " 553";
        when 552 => reg2_string <= " 552";
        when 551 => reg2_string <= " 551";
        when 550 => reg2_string <= " 550";
        when 549 => reg2_string <= " 549";
        when 548 => reg2_string <= " 548";
        when 547 => reg2_string <= " 547";
        when 546 => reg2_string <= " 546";
        when 545 => reg2_string <= " 545";
        when 544 => reg2_string <= " 544";
        when 543 => reg2_string <= " 543";
        when 542 => reg2_string <= " 542";
        when 541 => reg2_string <= " 541";
        when 540 => reg2_string <= " 540";
        when 539 => reg2_string <= " 539";
        when 538 => reg2_string <= " 538";
        when 537 => reg2_string <= " 537";
        when 536 => reg2_string <= " 536";
        when 535 => reg2_string <= " 535";
        when 534 => reg2_string <= " 534";
        when 533 => reg2_string <= " 533";
        when 532 => reg2_string <= " 532";
        when 531 => reg2_string <= " 531";
        when 530 => reg2_string <= " 530";
        when 529 => reg2_string <= " 529";
        when 528 => reg2_string <= " 528";
        when 527 => reg2_string <= " 527";
        when 526 => reg2_string <= " 526";
        when 525 => reg2_string <= " 525";
        when 524 => reg2_string <= " 524";
        when 523 => reg2_string <= " 523";
        when 522 => reg2_string <= " 522";
        when 521 => reg2_string <= " 521";
        when 520 => reg2_string <= " 520";
        when 519 => reg2_string <= " 519";
        when 518 => reg2_string <= " 518";
        when 517 => reg2_string <= " 517";
        when 516 => reg2_string <= " 516";
        when 515 => reg2_string <= " 515";
        when 514 => reg2_string <= " 514";
        when 513 => reg2_string <= " 513";
        when 512 => reg2_string <= " 512";
        when 511 => reg2_string <= " 511";
        when 510 => reg2_string <= " 510";
        when 509 => reg2_string <= " 509";
        when 508 => reg2_string <= " 508";
        when 507 => reg2_string <= " 507";
        when 506 => reg2_string <= " 506";
        when 505 => reg2_string <= " 505";
        when 504 => reg2_string <= " 504";
        when 503 => reg2_string <= " 503";
        when 502 => reg2_string <= " 502";
        when 501 => reg2_string <= " 501";
        when 500 => reg2_string <= " 500";
        when 499 => reg2_string <= " 499";
        when 498 => reg2_string <= " 498";
        when 497 => reg2_string <= " 497";
        when 496 => reg2_string <= " 496";
        when 495 => reg2_string <= " 495";
        when 494 => reg2_string <= " 494";
        when 493 => reg2_string <= " 493";
        when 492 => reg2_string <= " 492";
        when 491 => reg2_string <= " 491";
        when 490 => reg2_string <= " 490";
        when 489 => reg2_string <= " 489";
        when 488 => reg2_string <= " 488";
        when 487 => reg2_string <= " 487";
        when 486 => reg2_string <= " 486";
        when 485 => reg2_string <= " 485";
        when 484 => reg2_string <= " 484";
        when 483 => reg2_string <= " 483";
        when 482 => reg2_string <= " 482";
        when 481 => reg2_string <= " 481";
        when 480 => reg2_string <= " 480";
        when 479 => reg2_string <= " 479";
        when 478 => reg2_string <= " 478";
        when 477 => reg2_string <= " 477";
        when 476 => reg2_string <= " 476";
        when 475 => reg2_string <= " 475";
        when 474 => reg2_string <= " 474";
        when 473 => reg2_string <= " 473";
        when 472 => reg2_string <= " 472";
        when 471 => reg2_string <= " 471";
        when 470 => reg2_string <= " 470";
        when 469 => reg2_string <= " 469";
        when 468 => reg2_string <= " 468";
        when 467 => reg2_string <= " 467";
        when 466 => reg2_string <= " 466";
        when 465 => reg2_string <= " 465";
        when 464 => reg2_string <= " 464";
        when 463 => reg2_string <= " 463";
        when 462 => reg2_string <= " 462";
        when 461 => reg2_string <= " 461";
        when 460 => reg2_string <= " 460";
        when 459 => reg2_string <= " 459";
        when 458 => reg2_string <= " 458";
        when 457 => reg2_string <= " 457";
        when 456 => reg2_string <= " 456";
        when 455 => reg2_string <= " 455";
        when 454 => reg2_string <= " 454";
        when 453 => reg2_string <= " 453";
        when 452 => reg2_string <= " 452";
        when 451 => reg2_string <= " 451";
        when 450 => reg2_string <= " 450";
        when 449 => reg2_string <= " 449";
        when 448 => reg2_string <= " 448";
        when 447 => reg2_string <= " 447";
        when 446 => reg2_string <= " 446";
        when 445 => reg2_string <= " 445";
        when 444 => reg2_string <= " 444";
        when 443 => reg2_string <= " 443";
        when 442 => reg2_string <= " 442";
        when 441 => reg2_string <= " 441";
        when 440 => reg2_string <= " 440";
        when 439 => reg2_string <= " 439";
        when 438 => reg2_string <= " 438";
        when 437 => reg2_string <= " 437";
        when 436 => reg2_string <= " 436";
        when 435 => reg2_string <= " 435";
        when 434 => reg2_string <= " 434";
        when 433 => reg2_string <= " 433";
        when 432 => reg2_string <= " 432";
        when 431 => reg2_string <= " 431";
        when 430 => reg2_string <= " 430";
        when 429 => reg2_string <= " 429";
        when 428 => reg2_string <= " 428";
        when 427 => reg2_string <= " 427";
        when 426 => reg2_string <= " 426";
        when 425 => reg2_string <= " 425";
        when 424 => reg2_string <= " 424";
        when 423 => reg2_string <= " 423";
        when 422 => reg2_string <= " 422";
        when 421 => reg2_string <= " 421";
        when 420 => reg2_string <= " 420";
        when 419 => reg2_string <= " 419";
        when 418 => reg2_string <= " 418";
        when 417 => reg2_string <= " 417";
        when 416 => reg2_string <= " 416";
        when 415 => reg2_string <= " 415";
        when 414 => reg2_string <= " 414";
        when 413 => reg2_string <= " 413";
        when 412 => reg2_string <= " 412";
        when 411 => reg2_string <= " 411";
        when 410 => reg2_string <= " 410";
        when 409 => reg2_string <= " 409";
        when 408 => reg2_string <= " 408";
        when 407 => reg2_string <= " 407";
        when 406 => reg2_string <= " 406";
        when 405 => reg2_string <= " 405";
        when 404 => reg2_string <= " 404";
        when 403 => reg2_string <= " 403";
        when 402 => reg2_string <= " 402";
        when 401 => reg2_string <= " 401";
        when 400 => reg2_string <= " 400";
        when 399 => reg2_string <= " 399";
        when 398 => reg2_string <= " 398";
        when 397 => reg2_string <= " 397";
        when 396 => reg2_string <= " 396";
        when 395 => reg2_string <= " 395";
        when 394 => reg2_string <= " 394";
        when 393 => reg2_string <= " 393";
        when 392 => reg2_string <= " 392";
        when 391 => reg2_string <= " 391";
        when 390 => reg2_string <= " 390";
        when 389 => reg2_string <= " 389";
        when 388 => reg2_string <= " 388";
        when 387 => reg2_string <= " 387";
        when 386 => reg2_string <= " 386";
        when 385 => reg2_string <= " 385";
        when 384 => reg2_string <= " 384";
        when 383 => reg2_string <= " 383";
        when 382 => reg2_string <= " 382";
        when 381 => reg2_string <= " 381";
        when 380 => reg2_string <= " 380";
        when 379 => reg2_string <= " 379";
        when 378 => reg2_string <= " 378";
        when 377 => reg2_string <= " 377";
        when 376 => reg2_string <= " 376";
        when 375 => reg2_string <= " 375";
        when 374 => reg2_string <= " 374";
        when 373 => reg2_string <= " 373";
        when 372 => reg2_string <= " 372";
        when 371 => reg2_string <= " 371";
        when 370 => reg2_string <= " 370";
        when 369 => reg2_string <= " 369";
        when 368 => reg2_string <= " 368";
        when 367 => reg2_string <= " 367";
        when 366 => reg2_string <= " 366";
        when 365 => reg2_string <= " 365";
        when 364 => reg2_string <= " 364";
        when 363 => reg2_string <= " 363";
        when 362 => reg2_string <= " 362";
        when 361 => reg2_string <= " 361";
        when 360 => reg2_string <= " 360";
        when 359 => reg2_string <= " 359";
        when 358 => reg2_string <= " 358";
        when 357 => reg2_string <= " 357";
        when 356 => reg2_string <= " 356";
        when 355 => reg2_string <= " 355";
        when 354 => reg2_string <= " 354";
        when 353 => reg2_string <= " 353";
        when 352 => reg2_string <= " 352";
        when 351 => reg2_string <= " 351";
        when 350 => reg2_string <= " 350";
        when 349 => reg2_string <= " 349";
        when 348 => reg2_string <= " 348";
        when 347 => reg2_string <= " 347";
        when 346 => reg2_string <= " 346";
        when 345 => reg2_string <= " 345";
        when 344 => reg2_string <= " 344";
        when 343 => reg2_string <= " 343";
        when 342 => reg2_string <= " 342";
        when 341 => reg2_string <= " 341";
        when 340 => reg2_string <= " 340";
        when 339 => reg2_string <= " 339";
        when 338 => reg2_string <= " 338";
        when 337 => reg2_string <= " 337";
        when 336 => reg2_string <= " 336";
        when 335 => reg2_string <= " 335";
        when 334 => reg2_string <= " 334";
        when 333 => reg2_string <= " 333";
        when 332 => reg2_string <= " 332";
        when 331 => reg2_string <= " 331";
        when 330 => reg2_string <= " 330";
        when 329 => reg2_string <= " 329";
        when 328 => reg2_string <= " 328";
        when 327 => reg2_string <= " 327";
        when 326 => reg2_string <= " 326";
        when 325 => reg2_string <= " 325";
        when 324 => reg2_string <= " 324";
        when 323 => reg2_string <= " 323";
        when 322 => reg2_string <= " 322";
        when 321 => reg2_string <= " 321";
        when 320 => reg2_string <= " 320";
        when 319 => reg2_string <= " 319";
        when 318 => reg2_string <= " 318";
        when 317 => reg2_string <= " 317";
        when 316 => reg2_string <= " 316";
        when 315 => reg2_string <= " 315";
        when 314 => reg2_string <= " 314";
        when 313 => reg2_string <= " 313";
        when 312 => reg2_string <= " 312";
        when 311 => reg2_string <= " 311";
        when 310 => reg2_string <= " 310";
        when 309 => reg2_string <= " 309";
        when 308 => reg2_string <= " 308";
        when 307 => reg2_string <= " 307";
        when 306 => reg2_string <= " 306";
        when 305 => reg2_string <= " 305";
        when 304 => reg2_string <= " 304";
        when 303 => reg2_string <= " 303";
        when 302 => reg2_string <= " 302";
        when 301 => reg2_string <= " 301";
        when 300 => reg2_string <= " 300";
        when 299 => reg2_string <= " 299";
        when 298 => reg2_string <= " 298";
        when 297 => reg2_string <= " 297";
        when 296 => reg2_string <= " 296";
        when 295 => reg2_string <= " 295";
        when 294 => reg2_string <= " 294";
        when 293 => reg2_string <= " 293";
        when 292 => reg2_string <= " 292";
        when 291 => reg2_string <= " 291";
        when 290 => reg2_string <= " 290";
        when 289 => reg2_string <= " 289";
        when 288 => reg2_string <= " 288";
        when 287 => reg2_string <= " 287";
        when 286 => reg2_string <= " 286";
        when 285 => reg2_string <= " 285";
        when 284 => reg2_string <= " 284";
        when 283 => reg2_string <= " 283";
        when 282 => reg2_string <= " 282";
        when 281 => reg2_string <= " 281";
        when 280 => reg2_string <= " 280";
        when 279 => reg2_string <= " 279";
        when 278 => reg2_string <= " 278";
        when 277 => reg2_string <= " 277";
        when 276 => reg2_string <= " 276";
        when 275 => reg2_string <= " 275";
        when 274 => reg2_string <= " 274";
        when 273 => reg2_string <= " 273";
        when 272 => reg2_string <= " 272";
        when 271 => reg2_string <= " 271";
        when 270 => reg2_string <= " 270";
        when 269 => reg2_string <= " 269";
        when 268 => reg2_string <= " 268";
        when 267 => reg2_string <= " 267";
        when 266 => reg2_string <= " 266";
        when 265 => reg2_string <= " 265";
        when 264 => reg2_string <= " 264";
        when 263 => reg2_string <= " 263";
        when 262 => reg2_string <= " 262";
        when 261 => reg2_string <= " 261";
        when 260 => reg2_string <= " 260";
        when 259 => reg2_string <= " 259";
        when 258 => reg2_string <= " 258";
        when 257 => reg2_string <= " 257";
        when 256 => reg2_string <= " 256";
        when 255 => reg2_string <= " 255";
        when 254 => reg2_string <= " 254";
        when 253 => reg2_string <= " 253";
        when 252 => reg2_string <= " 252";
        when 251 => reg2_string <= " 251";
        when 250 => reg2_string <= " 250";
        when 249 => reg2_string <= " 249";
        when 248 => reg2_string <= " 248";
        when 247 => reg2_string <= " 247";
        when 246 => reg2_string <= " 246";
        when 245 => reg2_string <= " 245";
        when 244 => reg2_string <= " 244";
        when 243 => reg2_string <= " 243";
        when 242 => reg2_string <= " 242";
        when 241 => reg2_string <= " 241";
        when 240 => reg2_string <= " 240";
        when 239 => reg2_string <= " 239";
        when 238 => reg2_string <= " 238";
        when 237 => reg2_string <= " 237";
        when 236 => reg2_string <= " 236";
        when 235 => reg2_string <= " 235";
        when 234 => reg2_string <= " 234";
        when 233 => reg2_string <= " 233";
        when 232 => reg2_string <= " 232";
        when 231 => reg2_string <= " 231";
        when 230 => reg2_string <= " 230";
        when 229 => reg2_string <= " 229";
        when 228 => reg2_string <= " 228";
        when 227 => reg2_string <= " 227";
        when 226 => reg2_string <= " 226";
        when 225 => reg2_string <= " 225";
        when 224 => reg2_string <= " 224";
        when 223 => reg2_string <= " 223";
        when 222 => reg2_string <= " 222";
        when 221 => reg2_string <= " 221";
        when 220 => reg2_string <= " 220";
        when 219 => reg2_string <= " 219";
        when 218 => reg2_string <= " 218";
        when 217 => reg2_string <= " 217";
        when 216 => reg2_string <= " 216";
        when 215 => reg2_string <= " 215";
        when 214 => reg2_string <= " 214";
        when 213 => reg2_string <= " 213";
        when 212 => reg2_string <= " 212";
        when 211 => reg2_string <= " 211";
        when 210 => reg2_string <= " 210";
        when 209 => reg2_string <= " 209";
        when 208 => reg2_string <= " 208";
        when 207 => reg2_string <= " 207";
        when 206 => reg2_string <= " 206";
        when 205 => reg2_string <= " 205";
        when 204 => reg2_string <= " 204";
        when 203 => reg2_string <= " 203";
        when 202 => reg2_string <= " 202";
        when 201 => reg2_string <= " 201";
        when 200 => reg2_string <= " 200";
        when 199 => reg2_string <= " 199";
        when 198 => reg2_string <= " 198";
        when 197 => reg2_string <= " 197";
        when 196 => reg2_string <= " 196";
        when 195 => reg2_string <= " 195";
        when 194 => reg2_string <= " 194";
        when 193 => reg2_string <= " 193";
        when 192 => reg2_string <= " 192";
        when 191 => reg2_string <= " 191";
        when 190 => reg2_string <= " 190";
        when 189 => reg2_string <= " 189";
        when 188 => reg2_string <= " 188";
        when 187 => reg2_string <= " 187";
        when 186 => reg2_string <= " 186";
        when 185 => reg2_string <= " 185";
        when 184 => reg2_string <= " 184";
        when 183 => reg2_string <= " 183";
        when 182 => reg2_string <= " 182";
        when 181 => reg2_string <= " 181";
        when 180 => reg2_string <= " 180";
        when 179 => reg2_string <= " 179";
        when 178 => reg2_string <= " 178";
        when 177 => reg2_string <= " 177";
        when 176 => reg2_string <= " 176";
        when 175 => reg2_string <= " 175";
        when 174 => reg2_string <= " 174";
        when 173 => reg2_string <= " 173";
        when 172 => reg2_string <= " 172";
        when 171 => reg2_string <= " 171";
        when 170 => reg2_string <= " 170";
        when 169 => reg2_string <= " 169";
        when 168 => reg2_string <= " 168";
        when 167 => reg2_string <= " 167";
        when 166 => reg2_string <= " 166";
        when 165 => reg2_string <= " 165";
        when 164 => reg2_string <= " 164";
        when 163 => reg2_string <= " 163";
        when 162 => reg2_string <= " 162";
        when 161 => reg2_string <= " 161";
        when 160 => reg2_string <= " 160";
        when 159 => reg2_string <= " 159";
        when 158 => reg2_string <= " 158";
        when 157 => reg2_string <= " 157";
        when 156 => reg2_string <= " 156";
        when 155 => reg2_string <= " 155";
        when 154 => reg2_string <= " 154";
        when 153 => reg2_string <= " 153";
        when 152 => reg2_string <= " 152";
        when 151 => reg2_string <= " 151";
        when 150 => reg2_string <= " 150";
        when 149 => reg2_string <= " 149";
        when 148 => reg2_string <= " 148";
        when 147 => reg2_string <= " 147";
        when 146 => reg2_string <= " 146";
        when 145 => reg2_string <= " 145";
        when 144 => reg2_string <= " 144";
        when 143 => reg2_string <= " 143";
        when 142 => reg2_string <= " 142";
        when 141 => reg2_string <= " 141";
        when 140 => reg2_string <= " 140";
        when 139 => reg2_string <= " 139";
        when 138 => reg2_string <= " 138";
        when 137 => reg2_string <= " 137";
        when 136 => reg2_string <= " 136";
        when 135 => reg2_string <= " 135";
        when 134 => reg2_string <= " 134";
        when 133 => reg2_string <= " 133";
        when 132 => reg2_string <= " 132";
        when 131 => reg2_string <= " 131";
        when 130 => reg2_string <= " 130";
        when 129 => reg2_string <= " 129";
        when 128 => reg2_string <= " 128";
        when 127 => reg2_string <= " 127";
        when 126 => reg2_string <= " 126";
        when 125 => reg2_string <= " 125";
        when 124 => reg2_string <= " 124";
        when 123 => reg2_string <= " 123";
        when 122 => reg2_string <= " 122";
        when 121 => reg2_string <= " 121";
        when 120 => reg2_string <= " 120";
        when 119 => reg2_string <= " 119";
        when 118 => reg2_string <= " 118";
        when 117 => reg2_string <= " 117";
        when 116 => reg2_string <= " 116";
        when 115 => reg2_string <= " 115";
        when 114 => reg2_string <= " 114";
        when 113 => reg2_string <= " 113";
        when 112 => reg2_string <= " 112";
        when 111 => reg2_string <= " 111";
        when 110 => reg2_string <= " 110";
        when 109 => reg2_string <= " 109";
        when 108 => reg2_string <= " 108";
            when 107 => reg2_string <= " 107";                                                                                        
            when 106 => reg2_string <= " 106";                                                                                        
            when 105 => reg2_string <= " 105";                                                                                        
            when 104 => reg2_string <= " 104";                                                                                        
            when 103 => reg2_string <= " 103";                                                                                        
            when 102 => reg2_string <= " 102";                                                                                        
            when 101 => reg2_string <= " 101";                                                                                        
            when 100 => reg2_string <= " 100";                                                                                        
            when 99 => reg2_string <= "  99";                                                                                         
            when 98 => reg2_string <= "  98";                                                                                         
            when 97 => reg2_string <= "  97";                                                                                         
            when 96 => reg2_string <= "  96";                                                                                         
            when 95 => reg2_string <= "  95";                                                                                         
            when 94 => reg2_string <= "  94";                                                                                         
            when 93 => reg2_string <= "  93";                                                                                         
            when 92 => reg2_string <= "  92";                                                                                         
            when 91 => reg2_string <= "  91";                                                                                         
            when 90 => reg2_string <= "  90";                                                                                         
            when 89 => reg2_string <= "  89";                                                                                         
            when 88 => reg2_string <= "  88";                                                                                         
            when 87 => reg2_string <= "  87";                                                                                         
            when 86 => reg2_string <= "  86";                                                                                         
            when 85 => reg2_string <= "  85";                                                                                         
            when 84 => reg2_string <= "  84";                                                                                         
            when 83 => reg2_string <= "  83";                                                                                         
            when 82 => reg2_string <= "  82";                                                                                         
            when 81 => reg2_string <= "  81";                                                                                         
            when 80 => reg2_string <= "  80";                                                                                         
            when 79 => reg2_string <= "  79";                                                                                         
            when 78 => reg2_string <= "  78";                                                                                         
            when 77 => reg2_string <= "  77";
            when 76 => reg2_string <= "  76";                                                                                         
            when 75 => reg2_string <= "  75";                                                                                         
            when 74 => reg2_string <= "  74";                                                                                         
            when 73 => reg2_string <= "  73";                                                                                         
            when 72 => reg2_string <= "  72";                                                                                         
            when 71 => reg2_string <= "  71";                                                                                         
            when 70 => reg2_string <= "  70";                                                                                         
            when 69 => reg2_string <= "  69";                                                                                         
            when 68 => reg2_string <= "  68";                                                                                         
            when 67 => reg2_string <= "  67";                                                                                         
            when 66 => reg2_string <= "  66";                                                                                         
            when 65 => reg2_string <= "  65";                                                                                         
            when 64 => reg2_string <= "  64";                                                                                         
            when 63 => reg2_string <= "  63";                                                                                         
            when 62 => reg2_string <= "  62";                                                                                         
            when 61 => reg2_string <= "  61";                                                                                         
            when 60 => reg2_string <= "  60";                                                                                         
            when 59 => reg2_string <= "  59";                                                                                         
            when 58 => reg2_string <= "  58";                                                                                         
            when 57 => reg2_string <= "  57";                                                                                         
            when 56 => reg2_string <= "  56";                                                                                         
            when 55 => reg2_string <= "  55";                                                                                         
            when 54 => reg2_string <= "  54";                                                                                         
            when 53 => reg2_string <= "  53";                                                                                         
            when 52 => reg2_string <= "  52";                                                                                         
            when 51 => reg2_string <= "  51";                                                                                         
            when 50 => reg2_string <= "  50";                                                                                         
            when 49 => reg2_string <= "  49";                                                                                         
            when 48 => reg2_string <= "  48";                                                                                         
            when 47 => reg2_string <= "  47";
            when 46 => reg2_string <= "  46";                                                                                         
            when 45 => reg2_string <= "  45";                                                                                         
            when 44 => reg2_string <= "  44";                                                                                         
            when 43 => reg2_string <= "  43";                                                                                         
            when 42 => reg2_string <= "  42";                                                                                         
            when 41 => reg2_string <= "  41";                                                                                         
            when 40 => reg2_string <= "  40";                                                                                         
            when 39 => reg2_string <= "  39";                                                                                         
            when 38 => reg2_string <= "  38";                                                                                         
            when 37 => reg2_string <= "  37";                                                                                         
            when 36 => reg2_string <= "  36";                                                                                         
            when 35 => reg2_string <= "  35";                                                                                         
            when 34 => reg2_string <= "  34";                                                                                         
            when 33 => reg2_string <= "  33";                                                                                         
            when 32 => reg2_string <= "  32";                                                                                         
            when 31 => reg2_string <= "  31";                                                                                         
            when 30 => reg2_string <= "  30";                                                                                         
            when 29 => reg2_string <= "  29";                                                                                         
            when 28 => reg2_string <= "  28";                                                                                         
            when 27 => reg2_string <= "  27";                                                                                         
            when 26 => reg2_string <= "  26";                                                                                         
            when 25 => reg2_string <= "  25";                                                                                         
            when 24 => reg2_string <= "  24";                                                                                         
            when 23 => reg2_string <= "  23";
            when 22 => reg2_string <= "  22";                                                                                         
            when 21 => reg2_string <= "  21";                                                                                         
            when 20 => reg2_string <= "  20";                                                                                         
            when 19 => reg2_string <= "  19";                                                                                         
            when 18 => reg2_string <= "  18";                                                                                         
            when 17 => reg2_string <= "  17";                                                                                         
            when 16 => reg2_string <= "  16";                                                                                         
            when 15 => reg2_string <= "  15";                                                                                         
            when 14 => reg2_string <= "  14";                                                                                         
            when 13 => reg2_string <= "  13";                                                                                         
            when 12 => reg2_string <= "  12";                                                                                         
            when 11 => reg2_string <= "  11";                                                                                         
            when 10 => reg2_string <= "  10";                                                                                         
            when 9  => reg2_string <= "   9";                                                                                          
            when 8  => reg2_string <= "   8";                                                                                          
            when 7  => reg2_string <= "   7";                                                                                          
            when 6  => reg2_string <= "   6";                                                                                          
            when 5  => reg2_string <= "   5";                                                                                          
            when 4  => reg2_string <= "   4";                                                                                          
            when 3  => reg2_string <= "   3";                                                                                          
            when 2  => reg2_string <= "   2";                                                                                          
            when 1  => reg2_string <= "   1";                                                                                          
            when 0  => reg2_string <= "   0";
            when -1 => reg2_string <= "  -1";
            when -2 => reg2_string <= "  -2";
            when -3 => reg2_string <= "  -3";
            when -4 => reg2_string <= "  -4";
            when -5 => reg2_string <= "  -5";
            when -6 => reg2_string <= "  -6";
            when -7 => reg2_string <= "  -7";
            when -8 => reg2_string <= "  -8";
            when -9 => reg2_string <= "  -9";
            when -10 => reg2_string <= " -10";
            when -11 => reg2_string <= " -11";
            when -12 => reg2_string <= " -12";
            when -13 => reg2_string <= " -13";
            when -14 => reg2_string <= " -14";
            when -15 => reg2_string <= " -15";
            when -16 => reg2_string <= " -16";
            when -17 => reg2_string <= " -17";
            when -18 => reg2_string <= " -18";
            when -19 => reg2_string <= " -19";
            when -20 => reg2_string <= " -20";
            when -21 => reg2_string <= " -21";
            when -22 => reg2_string <= " -22";
            when -23 => reg2_string <= " -23";
            when -24 => reg2_string <= " -24";
            when -25 => reg2_string <= " -25";
            when -26 => reg2_string <= " -26";
            when -27 => reg2_string <= " -27";
            when -28 => reg2_string <= " -28";
            when -29 => reg2_string <= " -29";
            when -30 => reg2_string <= " -30";
            when -31 => reg2_string <= " -31";
            when -32 => reg2_string <= " -32";
            when -33 => reg2_string <= " -33";
            when -34 => reg2_string <= " -34";
            when -35 => reg2_string <= " -35";
            when -36 => reg2_string <= " -36";
            when -37 => reg2_string <= " -37";
            when -38 => reg2_string <= " -38";
            when -39 => reg2_string <= " -39";
            when -40 => reg2_string <= " -40";
            when -41 => reg2_string <= " -41";
            when -42 => reg2_string <= " -42";
            when -43 => reg2_string <= " -43";
            when -44 => reg2_string <= " -44";
            when -45 => reg2_string <= " -45";
            when -46 => reg2_string <= " -46";
            when -47 => reg2_string <= " -47";
            when -48 => reg2_string <= " -48";
            when -49 => reg2_string <= " -49";
            when -50 => reg2_string <= " -50";
            when -51 => reg2_string <= " -51";
            when -52 => reg2_string <= " -52";
            when -53 => reg2_string <= " -53";
            when -54 => reg2_string <= " -54";
            when -55 => reg2_string <= " -55";
            when -56 => reg2_string <= " -56";
            when -57 => reg2_string <= " -57";
            when -58 => reg2_string <= " -58";
            when -59 => reg2_string <= " -59";
            when -60 => reg2_string <= " -60";
            when -61 => reg2_string <= " -61";
            when -62 => reg2_string <= " -62";
            when -63 => reg2_string <= " -63";
            when -64 => reg2_string <= " -64";
            when -65 => reg2_string <= " -65";
            when -66 => reg2_string <= " -66";
            when -67 => reg2_string <= " -67";
            when -68 => reg2_string <= " -68";
            when -69 => reg2_string <= " -69";
            when -70 => reg2_string <= " -70";
            when -71 => reg2_string <= " -71";
            when -72 => reg2_string <= " -72";
            when -73 => reg2_string <= " -73";
            when -74 => reg2_string <= " -74";
            when -75 => reg2_string <= " -75";
            when -76 => reg2_string <= " -76";
            when -77 => reg2_string <= " -77";
            when -78 => reg2_string <= " -78";
            when -79 => reg2_string <= " -79";
            when -80 => reg2_string <= " -80";
            when -81 => reg2_string <= " -81";
            when -82 => reg2_string <= " -82";
            when -83 => reg2_string <= " -83";
            when -84 => reg2_string <= " -84";
            when -85 => reg2_string <= " -85";
            when -86 => reg2_string <= " -86";
            when -87 => reg2_string <= " -87";
            when -88 => reg2_string <= " -88";
            when -89 => reg2_string <= " -89";
            when -90 => reg2_string <= " -90";
            when -91 => reg2_string <= " -91";
            when -92 => reg2_string <= " -92";
            when -93 => reg2_string <= " -93";
            when -94 => reg2_string <= " -94";
            when -95 => reg2_string <= " -95";
            when -96 => reg2_string <= " -96";
            when -97 => reg2_string <= " -97";
            when -98 => reg2_string <= " -98";
            when -99 => reg2_string <= " -99";
            when -100 => reg2_string <= "-100";
            when -101 => reg2_string <= "-101";
            when -102 => reg2_string <= "-102";
            when -103 => reg2_string <= "-103";
            when -104 => reg2_string <= "-104";
            when -105 => reg2_string <= "-105";
            when -106 => reg2_string <= "-106";
            when -107 => reg2_string <= "-107";
            when -108 => reg2_string <= "-108";
            when -109 => reg2_string <= "-109";
            when -110 => reg2_string <= "-110";
            when -111 => reg2_string <= "-111";
            when -112 => reg2_string <= "-112";
            when -113 => reg2_string <= "-113";
            when -114 => reg2_string <= "-114";
            when -115 => reg2_string <= "-115";
            when -116 => reg2_string <= "-116";
            when -117 => reg2_string <= "-117";
            when -118 => reg2_string <= "-118";
            when -119 => reg2_string <= "-119";
            when -120 => reg2_string <= "-120";
            when -121 => reg2_string <= "-121";
            when -122 => reg2_string <= "-122";
            when -123 => reg2_string <= "-123";
            when -124 => reg2_string <= "-124";
            when -125 => reg2_string <= "-125";
            when -126 => reg2_string <= "-126";
            when -127 => reg2_string <= "-127";
            when -128 => reg2_string <= "-128";
            when -129 => reg2_string <= "-129";
            when -130 => reg2_string <= "-130";
            when -131 => reg2_string <= "-131";
            when -132 => reg2_string <= "-132";
            when -133 => reg2_string <= "-133";
            when -134 => reg2_string <= "-134";
            when -135 => reg2_string <= "-135";
            when -136 => reg2_string <= "-136";
            when -137 => reg2_string <= "-137";
            when -138 => reg2_string <= "-138";
            when -139 => reg2_string <= "-139";
            when -140 => reg2_string <= "-140";
            when -141 => reg2_string <= "-141";
            when -142 => reg2_string <= "-142";
            when -143 => reg2_string <= "-143";
            when -144 => reg2_string <= "-144";
            when -145 => reg2_string <= "-145";
            when -146 => reg2_string <= "-146";
            when -147 => reg2_string <= "-147";
            when -148 => reg2_string <= "-148";
            when -149 => reg2_string <= "-149";
            when -150 => reg2_string <= "-150";
            when -151 => reg2_string <= "-151";
            when -152 => reg2_string <= "-152";
            when -153 => reg2_string <= "-153";
            when -154 => reg2_string <= "-154";
            when -155 => reg2_string <= "-155";
            when -156 => reg2_string <= "-156";
            when -157 => reg2_string <= "-157";
            when -158 => reg2_string <= "-158";
            when -159 => reg2_string <= "-159";
            when -160 => reg2_string <= "-160";
            when -161 => reg2_string <= "-161";
            when -162 => reg2_string <= "-162";
            when -163 => reg2_string <= "-163";
            when -164 => reg2_string <= "-164";
            when -165 => reg2_string <= "-165";
            when -166 => reg2_string <= "-166";
            when -167 => reg2_string <= "-167";
            when -168 => reg2_string <= "-168";
            when -169 => reg2_string <= "-169";
            when -170 => reg2_string <= "-170";
            when -171 => reg2_string <= "-171";
            when -172 => reg2_string <= "-172";
            when -173 => reg2_string <= "-173";
            when -174 => reg2_string <= "-174";
            when -175 => reg2_string <= "-175";
            when -176 => reg2_string <= "-176";
            when -177 => reg2_string <= "-177";
            when -178 => reg2_string <= "-178";
            when -179 => reg2_string <= "-179";
            when -180 => reg2_string <= "-180";
            when -181 => reg2_string <= "-181";
            when -182 => reg2_string <= "-182";
            when -183 => reg2_string <= "-183";
            when -184 => reg2_string <= "-184";
            when -185 => reg2_string <= "-185";
            when -186 => reg2_string <= "-186";
            when -187 => reg2_string <= "-187";
            when -188 => reg2_string <= "-188";
            when -189 => reg2_string <= "-189";
            when -190 => reg2_string <= "-190";
            when -191 => reg2_string <= "-191";
            when -192 => reg2_string <= "-192";
            when -193 => reg2_string <= "-193";
            when -194 => reg2_string <= "-194";
            when -195 => reg2_string <= "-195";
            when -196 => reg2_string <= "-196";
            when -197 => reg2_string <= "-197";
            when -198 => reg2_string <= "-198";
            when -199 => reg2_string <= "-199";
            when -200 => reg2_string <= "-200";
            when -201 => reg2_string <= "-201";
            when -202 => reg2_string <= "-202";
            when -203 => reg2_string <= "-203";
            when -204 => reg2_string <= "-204";
            when -205 => reg2_string <= "-205";
            when -206 => reg2_string <= "-206";
            when -207 => reg2_string <= "-207";
            when -208 => reg2_string <= "-208";
            when -209 => reg2_string <= "-209";
            when -210 => reg2_string <= "-210";
            when -211 => reg2_string <= "-211";
            when -212 => reg2_string <= "-212";
            when -213 => reg2_string <= "-213";
            when -214 => reg2_string <= "-214";
            when -215 => reg2_string <= "-215";
            when -216 => reg2_string <= "-216";
            when -217 => reg2_string <= "-217";
            when -218 => reg2_string <= "-218";
            when -219 => reg2_string <= "-219";
            when -220 => reg2_string <= "-220";
            when -221 => reg2_string <= "-221";
            when -222 => reg2_string <= "-222";
            when -223 => reg2_string <= "-223";
            when -224 => reg2_string <= "-224";
            when -225 => reg2_string <= "-225";
            when -226 => reg2_string <= "-226";
            when -227 => reg2_string <= "-227";
            when -228 => reg2_string <= "-228";
            when -229 => reg2_string <= "-229";
            when -230 => reg2_string <= "-230";
            when -231 => reg2_string <= "-231";
            when -232 => reg2_string <= "-232";
            when -233 => reg2_string <= "-233";
            when -234 => reg2_string <= "-234";
            when -235 => reg2_string <= "-235";
            when -236 => reg2_string <= "-236";
            when -237 => reg2_string <= "-237";
            when -238 => reg2_string <= "-238";
            when -239 => reg2_string <= "-239";
            when -240 => reg2_string <= "-240";
            when -241 => reg2_string <= "-241";
            when -242 => reg2_string <= "-242";
            when -243 => reg2_string <= "-243";
            when -244 => reg2_string <= "-244";
            when -245 => reg2_string <= "-245";
            when -246 => reg2_string <= "-246";
            when -247 => reg2_string <= "-247";
            when -248 => reg2_string <= "-248";
            when -249 => reg2_string <= "-249";
            when -250 => reg2_string <= "-250";
            when -251 => reg2_string <= "-251";
            when -252 => reg2_string <= "-252";
            when -253 => reg2_string <= "-253";
            when -254 => reg2_string <= "-254";
            when -255 => reg2_string <= "-255";
            when -256 => reg2_string <= "-256";
            when -257 => reg2_string <= "-257";
            when -258 => reg2_string <= "-258";
            when -259 => reg2_string <= "-259";
            when -260 => reg2_string <= "-260";
            when -261 => reg2_string <= "-261";
            when -262 => reg2_string <= "-262";
            when -263 => reg2_string <= "-263";
            when -264 => reg2_string <= "-264";
            when -265 => reg2_string <= "-265";
            when -266 => reg2_string <= "-266";
            when -267 => reg2_string <= "-267";
            when -268 => reg2_string <= "-268";
            when -269 => reg2_string <= "-269";
            when -270 => reg2_string <= "-270";
            when -271 => reg2_string <= "-271";
            when -272 => reg2_string <= "-272";
            when -273 => reg2_string <= "-273";
            when -274 => reg2_string <= "-274";
            when -275 => reg2_string <= "-275";
            when -276 => reg2_string <= "-276";
            when -277 => reg2_string <= "-277";
            when -278 => reg2_string <= "-278";
            when -279 => reg2_string <= "-279";
            when -280 => reg2_string <= "-280";
            when -281 => reg2_string <= "-281";
            when -282 => reg2_string <= "-282";
            when -283 => reg2_string <= "-283";
            when -284 => reg2_string <= "-284";
            when -285 => reg2_string <= "-285";
            when -286 => reg2_string <= "-286";
            when -287 => reg2_string <= "-287";
            when -288 => reg2_string <= "-288";
            when -289 => reg2_string <= "-289";
            when -290 => reg2_string <= "-290";
            when -291 => reg2_string <= "-291";
            when -292 => reg2_string <= "-292";
            when -293 => reg2_string <= "-293";
            when -294 => reg2_string <= "-294";
            when -295 => reg2_string <= "-295";
            when -296 => reg2_string <= "-296";
            when -297 => reg2_string <= "-297";
            when -298 => reg2_string <= "-298";
            when -299 => reg2_string <= "-299";
            when -300 => reg2_string <= "-300";
            when -301 => reg2_string <= "-301";
            when -302 => reg2_string <= "-302";
            when -303 => reg2_string <= "-303";
            when -304 => reg2_string <= "-304";
            when -305 => reg2_string <= "-305";
            when -306 => reg2_string <= "-306";
            when -307 => reg2_string <= "-307";
            when -308 => reg2_string <= "-308";
            when -309 => reg2_string <= "-309";
            when -310 => reg2_string <= "-310";
            when -311 => reg2_string <= "-311";
            when -312 => reg2_string <= "-312";
            when -313 => reg2_string <= "-313";
            when -314 => reg2_string <= "-314";
            when -315 => reg2_string <= "-315";
            when -316 => reg2_string <= "-316";
            when -317 => reg2_string <= "-317";
            when -318 => reg2_string <= "-318";
            when -319 => reg2_string <= "-319";
            when -320 => reg2_string <= "-320";
            when -321 => reg2_string <= "-321";
            when -322 => reg2_string <= "-322";
            when -323 => reg2_string <= "-323";
            when -324 => reg2_string <= "-324";
            when -325 => reg2_string <= "-325";
            when -326 => reg2_string <= "-326";
            when -327 => reg2_string <= "-327";
            when -328 => reg2_string <= "-328";
            when -329 => reg2_string <= "-329";
            when -330 => reg2_string <= "-330";
            when -331 => reg2_string <= "-331";
            when -332 => reg2_string <= "-332";
            when -333 => reg2_string <= "-333";
            when -334 => reg2_string <= "-334";
            when -335 => reg2_string <= "-335";
            when -336 => reg2_string <= "-336";
            when -337 => reg2_string <= "-337";
            when -338 => reg2_string <= "-338";
            when -339 => reg2_string <= "-339";
            when -340 => reg2_string <= "-340";
            when -341 => reg2_string <= "-341";
            when -342 => reg2_string <= "-342";
            when -343 => reg2_string <= "-343";
            when -344 => reg2_string <= "-344";
            when -345 => reg2_string <= "-345";
            when -346 => reg2_string <= "-346";
            when -347 => reg2_string <= "-347";
            when -348 => reg2_string <= "-348";
            when -349 => reg2_string <= "-349";
            when -350 => reg2_string <= "-350";
            when -351 => reg2_string <= "-351";
            when -352 => reg2_string <= "-352";
            when -353 => reg2_string <= "-353";
            when -354 => reg2_string <= "-354";
            when -355 => reg2_string <= "-355";
            when -356 => reg2_string <= "-356";
            when -357 => reg2_string <= "-357";
            when -358 => reg2_string <= "-358";
            when -359 => reg2_string <= "-359";
            when -360 => reg2_string <= "-360";
            when -361 => reg2_string <= "-361";
            when -362 => reg2_string <= "-362";
            when -363 => reg2_string <= "-363";
            when -364 => reg2_string <= "-364";
            when -365 => reg2_string <= "-365";
            when -366 => reg2_string <= "-366";
            when -367 => reg2_string <= "-367";
            when -368 => reg2_string <= "-368";
            when -369 => reg2_string <= "-369";
            when -370 => reg2_string <= "-370";
            when -371 => reg2_string <= "-371";
            when -372 => reg2_string <= "-372";
            when -373 => reg2_string <= "-373";
            when -374 => reg2_string <= "-374";
            when -375 => reg2_string <= "-375";
            when -376 => reg2_string <= "-376";
            when -377 => reg2_string <= "-377";
            when -378 => reg2_string <= "-378";
            when -379 => reg2_string <= "-379";
            when -380 => reg2_string <= "-380";
            when -381 => reg2_string <= "-381";
            when -382 => reg2_string <= "-382";
            when -383 => reg2_string <= "-383";
            when -384 => reg2_string <= "-384";
            when -385 => reg2_string <= "-385";
            when -386 => reg2_string <= "-386";
            when -387 => reg2_string <= "-387";
            when -388 => reg2_string <= "-388";
            when -389 => reg2_string <= "-389";
            when -390 => reg2_string <= "-390";
            when -391 => reg2_string <= "-391";
            when -392 => reg2_string <= "-392";
            when -393 => reg2_string <= "-393";
            when -394 => reg2_string <= "-394";
            when -395 => reg2_string <= "-395";
            when -396 => reg2_string <= "-396";
            when -397 => reg2_string <= "-397";
            when -398 => reg2_string <= "-398";
            when -399 => reg2_string <= "-399";
            when -400 => reg2_string <= "-400";
            when -401 => reg2_string <= "-401";
            when -402 => reg2_string <= "-402";
            when -403 => reg2_string <= "-403";
            when -404 => reg2_string <= "-404";
            when -405 => reg2_string <= "-405";
            when -406 => reg2_string <= "-406";
            when -407 => reg2_string <= "-407";
            when -408 => reg2_string <= "-408";
            when -409 => reg2_string <= "-409";
            when -410 => reg2_string <= "-410";
            when -411 => reg2_string <= "-411";
            when -412 => reg2_string <= "-412";
            when -413 => reg2_string <= "-413";
            when -414 => reg2_string <= "-414";
            when -415 => reg2_string <= "-415";
            when -416 => reg2_string <= "-416";
            when -417 => reg2_string <= "-417";
            when -418 => reg2_string <= "-418";
            when -419 => reg2_string <= "-419";
            when -420 => reg2_string <= "-420";
            when -421 => reg2_string <= "-421";
            when -422 => reg2_string <= "-422";
            when -423 => reg2_string <= "-423";
            when -424 => reg2_string <= "-424";
            when -425 => reg2_string <= "-425";
            when -426 => reg2_string <= "-426";
            when -427 => reg2_string <= "-427";
            when -428 => reg2_string <= "-428";
            when -429 => reg2_string <= "-429";
            when -430 => reg2_string <= "-430";
            when -431 => reg2_string <= "-431";
            when -432 => reg2_string <= "-432";
            when -433 => reg2_string <= "-433";
            when -434 => reg2_string <= "-434";
            when -435 => reg2_string <= "-435";
            when -436 => reg2_string <= "-436";
            when -437 => reg2_string <= "-437";
            when -438 => reg2_string <= "-438";
            when -439 => reg2_string <= "-439";
            when -440 => reg2_string <= "-440";
            when -441 => reg2_string <= "-441";
            when -442 => reg2_string <= "-442";
            when -443 => reg2_string <= "-443";
            when -444 => reg2_string <= "-444";
            when -445 => reg2_string <= "-445";
            when -446 => reg2_string <= "-446";
            when -447 => reg2_string <= "-447";
            when -448 => reg2_string <= "-448";
            when -449 => reg2_string <= "-449";
            when -450 => reg2_string <= "-450";
            when -451 => reg2_string <= "-451";
            when -452 => reg2_string <= "-452";
            when -453 => reg2_string <= "-453";
            when -454 => reg2_string <= "-454";
            when -455 => reg2_string <= "-455";
            when -456 => reg2_string <= "-456";
            when -457 => reg2_string <= "-457";
            when -458 => reg2_string <= "-458";
            when -459 => reg2_string <= "-459";
            when -460 => reg2_string <= "-460";
            when -461 => reg2_string <= "-461";
            when -462 => reg2_string <= "-462";
            when -463 => reg2_string <= "-463";
            when -464 => reg2_string <= "-464";
            when -465 => reg2_string <= "-465";
            when -466 => reg2_string <= "-466";
            when -467 => reg2_string <= "-467";
            when -468 => reg2_string <= "-468";
            when -469 => reg2_string <= "-469";
            when -470 => reg2_string <= "-470";
            when -471 => reg2_string <= "-471";
            when -472 => reg2_string <= "-472";
            when -473 => reg2_string <= "-473";
            when -474 => reg2_string <= "-474";
            when -475 => reg2_string <= "-475";
            when -476 => reg2_string <= "-476";
            when -477 => reg2_string <= "-477";
            when -478 => reg2_string <= "-478";
            when -479 => reg2_string <= "-479";
            when -480 => reg2_string <= "-480";
            when -481 => reg2_string <= "-481";
            when -482 => reg2_string <= "-482";
            when -483 => reg2_string <= "-483";
            when -484 => reg2_string <= "-484";
            when -485 => reg2_string <= "-485";
            when -486 => reg2_string <= "-486";
            when -487 => reg2_string <= "-487";
            when -488 => reg2_string <= "-488";
            when -489 => reg2_string <= "-489";
            when -490 => reg2_string <= "-490";
            when -491 => reg2_string <= "-491";
            when -492 => reg2_string <= "-492";
            when -493 => reg2_string <= "-493";
            when -494 => reg2_string <= "-494";
            when -495 => reg2_string <= "-495";
            when -496 => reg2_string <= "-496";
            when -497 => reg2_string <= "-497";
            when -498 => reg2_string <= "-498";
            when -499 => reg2_string <= "-499";
            when -500 => reg2_string <= "-500";
            when -501 => reg2_string <= "-501";
            when -502 => reg2_string <= "-502";
            when -503 => reg2_string <= "-503";
            when -504 => reg2_string <= "-504";
            when -505 => reg2_string <= "-505";
            when -506 => reg2_string <= "-506";
            when -507 => reg2_string <= "-507";
            when -508 => reg2_string <= "-508";
            when -509 => reg2_string <= "-509";
            when -510 => reg2_string <= "-510";
            when -511 => reg2_string <= "-511";
            when -512 => reg2_string <= "-512";
            when -513 => reg2_string <= "-513";
            when -514 => reg2_string <= "-514";
            when -515 => reg2_string <= "-515";
            when -516 => reg2_string <= "-516";
            when -517 => reg2_string <= "-517";
            when -518 => reg2_string <= "-518";
            when -519 => reg2_string <= "-519";
            when -520 => reg2_string <= "-520";
            when -521 => reg2_string <= "-521";
            when -522 => reg2_string <= "-522";
            when -523 => reg2_string <= "-523";
            when -524 => reg2_string <= "-524";
            when -525 => reg2_string <= "-525";
            when -526 => reg2_string <= "-526";
            when -527 => reg2_string <= "-527";
            when -528 => reg2_string <= "-528";
            when -529 => reg2_string <= "-529";
            when -530 => reg2_string <= "-530";
            when -531 => reg2_string <= "-531";
            when -532 => reg2_string <= "-532";
            when -533 => reg2_string <= "-533";
            when -534 => reg2_string <= "-534";
            when -535 => reg2_string <= "-535";
            when -536 => reg2_string <= "-536";
            when -537 => reg2_string <= "-537";
            when -538 => reg2_string <= "-538";
            when -539 => reg2_string <= "-539";
            when -540 => reg2_string <= "-540";
            when -541 => reg2_string <= "-541";
            when -542 => reg2_string <= "-542";
            when -543 => reg2_string <= "-543";
            when -544 => reg2_string <= "-544";
            when -545 => reg2_string <= "-545";
            when -546 => reg2_string <= "-546";
            when -547 => reg2_string <= "-547";
            when -548 => reg2_string <= "-548";
            when -549 => reg2_string <= "-549";
            when -550 => reg2_string <= "-550";
            when -551 => reg2_string <= "-551";
            when -552 => reg2_string <= "-552";
            when -553 => reg2_string <= "-553";
            when -554 => reg2_string <= "-554";
            when -555 => reg2_string <= "-555";
            when -556 => reg2_string <= "-556";
            when -557 => reg2_string <= "-557";
            when -558 => reg2_string <= "-558";
            when -559 => reg2_string <= "-559";
            when -560 => reg2_string <= "-560";
            when -561 => reg2_string <= "-561";
            when -562 => reg2_string <= "-562";
            when -563 => reg2_string <= "-563";
            when -564 => reg2_string <= "-564";
            when -565 => reg2_string <= "-565";
            when -566 => reg2_string <= "-566";
            when -567 => reg2_string <= "-567";
            when -568 => reg2_string <= "-568";
            when -569 => reg2_string <= "-569";
            when -570 => reg2_string <= "-570";
            when -571 => reg2_string <= "-571";
            when -572 => reg2_string <= "-572";
            when -573 => reg2_string <= "-573";
            when -574 => reg2_string <= "-574";
            when -575 => reg2_string <= "-575";
            when -576 => reg2_string <= "-576";
            when -577 => reg2_string <= "-577";
            when -578 => reg2_string <= "-578";
            when -579 => reg2_string <= "-579";
            when -580 => reg2_string <= "-580";
            when -581 => reg2_string <= "-581";
            when -582 => reg2_string <= "-582";
            when -583 => reg2_string <= "-583";
            when -584 => reg2_string <= "-584";
            when -585 => reg2_string <= "-585";
            when -586 => reg2_string <= "-586";
            when -587 => reg2_string <= "-587";
            when -588 => reg2_string <= "-588";
            when -589 => reg2_string <= "-589";
            when -590 => reg2_string <= "-590";
            when -591 => reg2_string <= "-591";
            when -592 => reg2_string <= "-592";
            when -593 => reg2_string <= "-593";
            when -594 => reg2_string <= "-594";
            when -595 => reg2_string <= "-595";
            when -596 => reg2_string <= "-596";
            when -597 => reg2_string <= "-597";
            when -598 => reg2_string <= "-598";
            when -599 => reg2_string <= "-599";
            when -600 => reg2_string <= "-600";
            when -601 => reg2_string <= "-601";
            when -602 => reg2_string <= "-602";
            when -603 => reg2_string <= "-603";
            when -604 => reg2_string <= "-604";
            when -605 => reg2_string <= "-605";
            when -606 => reg2_string <= "-606";
            when -607 => reg2_string <= "-607";
            when -608 => reg2_string <= "-608";
            when -609 => reg2_string <= "-609";
            when -610 => reg2_string <= "-610";
            when -611 => reg2_string <= "-611";
            when -612 => reg2_string <= "-612";
            when -613 => reg2_string <= "-613";
            when -614 => reg2_string <= "-614";
            when -615 => reg2_string <= "-615";
            when -616 => reg2_string <= "-616";
            when -617 => reg2_string <= "-617";
            when -618 => reg2_string <= "-618";
            when -619 => reg2_string <= "-619";
            when -620 => reg2_string <= "-620";
            when -621 => reg2_string <= "-621";
            when -622 => reg2_string <= "-622";
            when -623 => reg2_string <= "-623";
            when -624 => reg2_string <= "-624";
            when -625 => reg2_string <= "-625";
            when -626 => reg2_string <= "-626";
            when -627 => reg2_string <= "-627";
            when -628 => reg2_string <= "-628";
            when -629 => reg2_string <= "-629";
            when -630 => reg2_string <= "-630";
            when -631 => reg2_string <= "-631";
            when -632 => reg2_string <= "-632";
            when -633 => reg2_string <= "-633";
            when -634 => reg2_string <= "-634";
            when -635 => reg2_string <= "-635";
            when -636 => reg2_string <= "-636";
            when -637 => reg2_string <= "-637";
            when -638 => reg2_string <= "-638";
            when -639 => reg2_string <= "-639";
            when -640 => reg2_string <= "-640";
            when -641 => reg2_string <= "-641";
            when -642 => reg2_string <= "-642";
            when -643 => reg2_string <= "-643";
            when -644 => reg2_string <= "-644";
            when -645 => reg2_string <= "-645";
            when -646 => reg2_string <= "-646";
            when -647 => reg2_string <= "-647";
            when -648 => reg2_string <= "-648";
            when -649 => reg2_string <= "-649";
            when -650 => reg2_string <= "-650";
            when -651 => reg2_string <= "-651";
            when -652 => reg2_string <= "-652";
            when -653 => reg2_string <= "-653";
            when -654 => reg2_string <= "-654";
            when -655 => reg2_string <= "-655";
            when -656 => reg2_string <= "-656";
            when -657 => reg2_string <= "-657";
            when -658 => reg2_string <= "-658";
            when -659 => reg2_string <= "-659";
            when -660 => reg2_string <= "-660";
            when -661 => reg2_string <= "-661";
            when -662 => reg2_string <= "-662";
            when -663 => reg2_string <= "-663";
            when -664 => reg2_string <= "-664";
            when -665 => reg2_string <= "-665";
            when -666 => reg2_string <= "-666";
            when -667 => reg2_string <= "-667";
            when -668 => reg2_string <= "-668";
            when -669 => reg2_string <= "-669";
            when -670 => reg2_string <= "-670";
            when -671 => reg2_string <= "-671";
            when -672 => reg2_string <= "-672";
            when -673 => reg2_string <= "-673";
            when -674 => reg2_string <= "-674";
            when -675 => reg2_string <= "-675";
            when -676 => reg2_string <= "-676";
            when -677 => reg2_string <= "-677";
            when -678 => reg2_string <= "-678";
            when -679 => reg2_string <= "-679";
            when -680 => reg2_string <= "-680";
            when -681 => reg2_string <= "-681";
            when -682 => reg2_string <= "-682";
            when -683 => reg2_string <= "-683";
            when -684 => reg2_string <= "-684";
            when -685 => reg2_string <= "-685";
            when -686 => reg2_string <= "-686";
            when -687 => reg2_string <= "-687";
            when -688 => reg2_string <= "-688";
            when -689 => reg2_string <= "-689";
            when -690 => reg2_string <= "-690";
            when -691 => reg2_string <= "-691";
            when -692 => reg2_string <= "-692";
            when -693 => reg2_string <= "-693";
            when -694 => reg2_string <= "-694";
            when -695 => reg2_string <= "-695";
            when -696 => reg2_string <= "-696";
            when -697 => reg2_string <= "-697";
            when -698 => reg2_string <= "-698";
            when -699 => reg2_string <= "-699";
            when -700 => reg2_string <= "-700";
            when -701 => reg2_string <= "-701";
            when -702 => reg2_string <= "-702";
            when -703 => reg2_string <= "-703";
            when -704 => reg2_string <= "-704";
            when -705 => reg2_string <= "-705";
            when -706 => reg2_string <= "-706";
            when -707 => reg2_string <= "-707";
            when -708 => reg2_string <= "-708";
            when -709 => reg2_string <= "-709";
            when -710 => reg2_string <= "-710";
            when -711 => reg2_string <= "-711";
            when -712 => reg2_string <= "-712";
            when -713 => reg2_string <= "-713";
            when -714 => reg2_string <= "-714";
            when -715 => reg2_string <= "-715";
            when -716 => reg2_string <= "-716";
            when -717 => reg2_string <= "-717";
            when -718 => reg2_string <= "-718";
            when -719 => reg2_string <= "-719";
            when -720 => reg2_string <= "-720";
            when -721 => reg2_string <= "-721";
            when -722 => reg2_string <= "-722";
            when -723 => reg2_string <= "-723";
            when -724 => reg2_string <= "-724";
            when -725 => reg2_string <= "-725";
            when -726 => reg2_string <= "-726";
            when -727 => reg2_string <= "-727";
            when -728 => reg2_string <= "-728";
            when -729 => reg2_string <= "-729";
            when -730 => reg2_string <= "-730";
            when -731 => reg2_string <= "-731";
            when -732 => reg2_string <= "-732";
            when -733 => reg2_string <= "-733";
            when -734 => reg2_string <= "-734";
            when -735 => reg2_string <= "-735";
            when -736 => reg2_string <= "-736";
            when -737 => reg2_string <= "-737";
            when -738 => reg2_string <= "-738";
            when -739 => reg2_string <= "-739";
            when -740 => reg2_string <= "-740";
            when -741 => reg2_string <= "-741";
            when -742 => reg2_string <= "-742";
            when -743 => reg2_string <= "-743";
            when -744 => reg2_string <= "-744";
            when -745 => reg2_string <= "-745";
            when -746 => reg2_string <= "-746";
            when -747 => reg2_string <= "-747";
            when -748 => reg2_string <= "-748";
            when -749 => reg2_string <= "-749";
            when -750 => reg2_string <= "-750";
            when -751 => reg2_string <= "-751";
            when -752 => reg2_string <= "-752";
            when -753 => reg2_string <= "-753";
            when -754 => reg2_string <= "-754";
            when -755 => reg2_string <= "-755";
            when -756 => reg2_string <= "-756";
            when -757 => reg2_string <= "-757";
            when -758 => reg2_string <= "-758";
            when -759 => reg2_string <= "-759";
            when -760 => reg2_string <= "-760";
            when -761 => reg2_string <= "-761";
            when -762 => reg2_string <= "-762";
            when -763 => reg2_string <= "-763";
            when -764 => reg2_string <= "-764";
            when -765 => reg2_string <= "-765";
            when -766 => reg2_string <= "-766";
            when -767 => reg2_string <= "-767";
            when -768 => reg2_string <= "-768";
            when -769 => reg2_string <= "-769";
            when -770 => reg2_string <= "-770";
            when -771 => reg2_string <= "-771";
            when -772 => reg2_string <= "-772";
            when -773 => reg2_string <= "-773";
            when -774 => reg2_string <= "-774";
            when -775 => reg2_string <= "-775";
            when -776 => reg2_string <= "-776";
            when -777 => reg2_string <= "-777";
            when -778 => reg2_string <= "-778";
            when -779 => reg2_string <= "-779";
            when -780 => reg2_string <= "-780";
            when -781 => reg2_string <= "-781";
            when -782 => reg2_string <= "-782";
            when -783 => reg2_string <= "-783";
            when -784 => reg2_string <= "-784";
            when -785 => reg2_string <= "-785";
            when -786 => reg2_string <= "-786";
            when -787 => reg2_string <= "-787";
            when -788 => reg2_string <= "-788";
            when -789 => reg2_string <= "-789";
            when -790 => reg2_string <= "-790";
            when -791 => reg2_string <= "-791";
            when -792 => reg2_string <= "-792";
            when -793 => reg2_string <= "-793";
            when -794 => reg2_string <= "-794";
            when -795 => reg2_string <= "-795";
            when -796 => reg2_string <= "-796";
            when -797 => reg2_string <= "-797";
            when -798 => reg2_string <= "-798";
            when -799 => reg2_string <= "-799";
            when -800 => reg2_string <= "-800";
            when -801 => reg2_string <= "-801";
            when -802 => reg2_string <= "-802";
            when -803 => reg2_string <= "-803";
            when -804 => reg2_string <= "-804";
            when -805 => reg2_string <= "-805";
            when -806 => reg2_string <= "-806";
            when -807 => reg2_string <= "-807";
            when -808 => reg2_string <= "-808";
            when -809 => reg2_string <= "-809";
            when -810 => reg2_string <= "-810";
            when -811 => reg2_string <= "-811";
            when -812 => reg2_string <= "-812";
            when -813 => reg2_string <= "-813";
            when -814 => reg2_string <= "-814";
            when -815 => reg2_string <= "-815";
            when -816 => reg2_string <= "-816";
            when -817 => reg2_string <= "-817";
            when -818 => reg2_string <= "-818";
            when -819 => reg2_string <= "-819";
            when -820 => reg2_string <= "-820";
            when -821 => reg2_string <= "-821";
            when -822 => reg2_string <= "-822";
            when -823 => reg2_string <= "-823";
            when -824 => reg2_string <= "-824";
            when -825 => reg2_string <= "-825";
            when -826 => reg2_string <= "-826";
            when -827 => reg2_string <= "-827";
            when -828 => reg2_string <= "-828";
            when -829 => reg2_string <= "-829";
            when -830 => reg2_string <= "-830";
            when -831 => reg2_string <= "-831";
            when -832 => reg2_string <= "-832";
            when -833 => reg2_string <= "-833";
            when -834 => reg2_string <= "-834";
            when -835 => reg2_string <= "-835";
            when -836 => reg2_string <= "-836";
            when -837 => reg2_string <= "-837";
            when -838 => reg2_string <= "-838";
            when -839 => reg2_string <= "-839";
            when -840 => reg2_string <= "-840";
            when -841 => reg2_string <= "-841";
            when -842 => reg2_string <= "-842";
            when -843 => reg2_string <= "-843";
            when -844 => reg2_string <= "-844";
            when -845 => reg2_string <= "-845";
            when -846 => reg2_string <= "-846";
            when -847 => reg2_string <= "-847";
            when -848 => reg2_string <= "-848";
            when -849 => reg2_string <= "-849";
            when -850 => reg2_string <= "-850";
            when -851 => reg2_string <= "-851";
            when -852 => reg2_string <= "-852";
            when -853 => reg2_string <= "-853";
            when -854 => reg2_string <= "-854";
            when -855 => reg2_string <= "-855";
            when -856 => reg2_string <= "-856";
            when -857 => reg2_string <= "-857";
            when -858 => reg2_string <= "-858";
            when -859 => reg2_string <= "-859";
            when -860 => reg2_string <= "-860";
            when -861 => reg2_string <= "-861";
            when -862 => reg2_string <= "-862";
            when -863 => reg2_string <= "-863";
            when -864 => reg2_string <= "-864";
            when -865 => reg2_string <= "-865";
            when -866 => reg2_string <= "-866";
            when -867 => reg2_string <= "-867";
            when -868 => reg2_string <= "-868";
            when -869 => reg2_string <= "-869";
            when -870 => reg2_string <= "-870";
            when -871 => reg2_string <= "-871";
            when -872 => reg2_string <= "-872";
            when -873 => reg2_string <= "-873";
            when -874 => reg2_string <= "-874";
            when -875 => reg2_string <= "-875";
            when -876 => reg2_string <= "-876";
            when -877 => reg2_string <= "-877";
            when -878 => reg2_string <= "-878";
            when -879 => reg2_string <= "-879";
            when -880 => reg2_string <= "-880";
            when -881 => reg2_string <= "-881";
            when -882 => reg2_string <= "-882";
            when -883 => reg2_string <= "-883";
            when -884 => reg2_string <= "-884";
            when -885 => reg2_string <= "-885";
            when -886 => reg2_string <= "-886";
            when -887 => reg2_string <= "-887";
            when -888 => reg2_string <= "-888";
            when -889 => reg2_string <= "-889";
            when -890 => reg2_string <= "-890";
            when -891 => reg2_string <= "-891";
            when -892 => reg2_string <= "-892";
            when -893 => reg2_string <= "-893";
            when -894 => reg2_string <= "-894";
            when -895 => reg2_string <= "-895";
            when -896 => reg2_string <= "-896";
            when -897 => reg2_string <= "-897";
            when -898 => reg2_string <= "-898";
            when -899 => reg2_string <= "-899";
            when -900 => reg2_string <= "-900";
            when -901 => reg2_string <= "-901";
            when -902 => reg2_string <= "-902";
            when -903 => reg2_string <= "-903";
            when -904 => reg2_string <= "-904";
            when -905 => reg2_string <= "-905";
            when -906 => reg2_string <= "-906";
            when -907 => reg2_string <= "-907";
            when -908 => reg2_string <= "-908";
            when -909 => reg2_string <= "-909";
            when -910 => reg2_string <= "-910";
            when -911 => reg2_string <= "-911";
            when -912 => reg2_string <= "-912";
            when -913 => reg2_string <= "-913";
            when -914 => reg2_string <= "-914";
            when -915 => reg2_string <= "-915";
            when -916 => reg2_string <= "-916";
            when -917 => reg2_string <= "-917";
            when -918 => reg2_string <= "-918";
            when -919 => reg2_string <= "-919";
            when -920 => reg2_string <= "-920";
            when -921 => reg2_string <= "-921";
            when -922 => reg2_string <= "-922";
            when -923 => reg2_string <= "-923";
            when -924 => reg2_string <= "-924";
            when -925 => reg2_string <= "-925";
            when -926 => reg2_string <= "-926";
            when -927 => reg2_string <= "-927";
            when -928 => reg2_string <= "-928";
            when -929 => reg2_string <= "-929";
            when -930 => reg2_string <= "-930";
            when -931 => reg2_string <= "-931";
            when -932 => reg2_string <= "-932";
            when -933 => reg2_string <= "-933";
            when -934 => reg2_string <= "-934";
            when -935 => reg2_string <= "-935";
            when -936 => reg2_string <= "-936";
            when -937 => reg2_string <= "-937";
            when -938 => reg2_string <= "-938";
            when -939 => reg2_string <= "-939";
            when -940 => reg2_string <= "-940";
            when -941 => reg2_string <= "-941";
            when -942 => reg2_string <= "-942";
            when -943 => reg2_string <= "-943";
            when -944 => reg2_string <= "-944";
            when -945 => reg2_string <= "-945";
            when -946 => reg2_string <= "-946";
            when -947 => reg2_string <= "-947";
            when -948 => reg2_string <= "-948";
            when -949 => reg2_string <= "-949";
            when -950 => reg2_string <= "-950";
            when -951 => reg2_string <= "-951";
            when -952 => reg2_string <= "-952";
            when -953 => reg2_string <= "-953";
            when -954 => reg2_string <= "-954";
            when -955 => reg2_string <= "-955";
            when -956 => reg2_string <= "-956";
            when -957 => reg2_string <= "-957";
            when -958 => reg2_string <= "-958";
            when -959 => reg2_string <= "-959";
            when -960 => reg2_string <= "-960";
            when -961 => reg2_string <= "-961";
            when -962 => reg2_string <= "-962";
            when -963 => reg2_string <= "-963";
            when -964 => reg2_string <= "-964";
            when -965 => reg2_string <= "-965";
            when -966 => reg2_string <= "-966";
            when -967 => reg2_string <= "-967";
            when -968 => reg2_string <= "-968";
            when -969 => reg2_string <= "-969";
            when -970 => reg2_string <= "-970";
            when -971 => reg2_string <= "-971";
            when -972 => reg2_string <= "-972";
            when -973 => reg2_string <= "-973";
            when -974 => reg2_string <= "-974";
            when -975 => reg2_string <= "-975";
            when -976 => reg2_string <= "-976";
            when -977 => reg2_string <= "-977";
            when -978 => reg2_string <= "-978";
            when -979 => reg2_string <= "-979";
            when -980 => reg2_string <= "-980";
            when -981 => reg2_string <= "-981";
            when -982 => reg2_string <= "-982";
            when -983 => reg2_string <= "-983";
            when -984 => reg2_string <= "-984";
            when -985 => reg2_string <= "-985";
            when -986 => reg2_string <= "-986";
            when -987 => reg2_string <= "-987";
            when -988 => reg2_string <= "-988";
            when -989 => reg2_string <= "-989";
            when -990 => reg2_string <= "-990";
            when -991 => reg2_string <= "-991";
            when -992 => reg2_string <= "-992";
            when -993 => reg2_string <= "-993";
            when -994 => reg2_string <= "-994";
            when -995 => reg2_string <= "-995";
            when -996 => reg2_string <= "-996";
            when -997 => reg2_string <= "-997";
            when -998 => reg2_string <= "-998";
            when -999 => reg2_string <= "-999";
            when others => reg2_string <= "    ";
        end case;
        
        case (reg1_int) is 
        when 999 => reg1_string <= " 999";
        when 998 => reg1_string <= " 998";
        when 997 => reg1_string <= " 997";
        when 996 => reg1_string <= " 996";
        when 995 => reg1_string <= " 995";
        when 994 => reg1_string <= " 994";
        when 993 => reg1_string <= " 993";
        when 992 => reg1_string <= " 992";
        when 991 => reg1_string <= " 991";
        when 990 => reg1_string <= " 990";
        when 989 => reg1_string <= " 989";
        when 988 => reg1_string <= " 988";
        when 987 => reg1_string <= " 987";
        when 986 => reg1_string <= " 986";
        when 985 => reg1_string <= " 985";
        when 984 => reg1_string <= " 984";
        when 983 => reg1_string <= " 983";
        when 982 => reg1_string <= " 982";
        when 981 => reg1_string <= " 981";
        when 980 => reg1_string <= " 980";
        when 979 => reg1_string <= " 979";
        when 978 => reg1_string <= " 978";
        when 977 => reg1_string <= " 977";
        when 976 => reg1_string <= " 976";
        when 975 => reg1_string <= " 975";
        when 974 => reg1_string <= " 974";
        when 973 => reg1_string <= " 973";
        when 972 => reg1_string <= " 972";
        when 971 => reg1_string <= " 971";
        when 970 => reg1_string <= " 970";
        when 969 => reg1_string <= " 969";
        when 968 => reg1_string <= " 968";
        when 967 => reg1_string <= " 967";
        when 966 => reg1_string <= " 966";
        when 965 => reg1_string <= " 965";
        when 964 => reg1_string <= " 964";
        when 963 => reg1_string <= " 963";
        when 962 => reg1_string <= " 962";
        when 961 => reg1_string <= " 961";
        when 960 => reg1_string <= " 960";
        when 959 => reg1_string <= " 959";
        when 958 => reg1_string <= " 958";
        when 957 => reg1_string <= " 957";
        when 956 => reg1_string <= " 956";
        when 955 => reg1_string <= " 955";
        when 954 => reg1_string <= " 954";
        when 953 => reg1_string <= " 953";
        when 952 => reg1_string <= " 952";
        when 951 => reg1_string <= " 951";
        when 950 => reg1_string <= " 950";
        when 949 => reg1_string <= " 949";
        when 948 => reg1_string <= " 948";
        when 947 => reg1_string <= " 947";
        when 946 => reg1_string <= " 946";
        when 945 => reg1_string <= " 945";
        when 944 => reg1_string <= " 944";
        when 943 => reg1_string <= " 943";
        when 942 => reg1_string <= " 942";
        when 941 => reg1_string <= " 941";
        when 940 => reg1_string <= " 940";
        when 939 => reg1_string <= " 939";
        when 938 => reg1_string <= " 938";
        when 937 => reg1_string <= " 937";
        when 936 => reg1_string <= " 936";
        when 935 => reg1_string <= " 935";
        when 934 => reg1_string <= " 934";
        when 933 => reg1_string <= " 933";
        when 932 => reg1_string <= " 932";
        when 931 => reg1_string <= " 931";
        when 930 => reg1_string <= " 930";
        when 929 => reg1_string <= " 929";
        when 928 => reg1_string <= " 928";
        when 927 => reg1_string <= " 927";
        when 926 => reg1_string <= " 926";
        when 925 => reg1_string <= " 925";
        when 924 => reg1_string <= " 924";
        when 923 => reg1_string <= " 923";
        when 922 => reg1_string <= " 922";
        when 921 => reg1_string <= " 921";
        when 920 => reg1_string <= " 920";
        when 919 => reg1_string <= " 919";
        when 918 => reg1_string <= " 918";
        when 917 => reg1_string <= " 917";
        when 916 => reg1_string <= " 916";
        when 915 => reg1_string <= " 915";
        when 914 => reg1_string <= " 914";
        when 913 => reg1_string <= " 913";
        when 912 => reg1_string <= " 912";
        when 911 => reg1_string <= " 911";
        when 910 => reg1_string <= " 910";
        when 909 => reg1_string <= " 909";
        when 908 => reg1_string <= " 908";
        when 907 => reg1_string <= " 907";
        when 906 => reg1_string <= " 906";
        when 905 => reg1_string <= " 905";
        when 904 => reg1_string <= " 904";
        when 903 => reg1_string <= " 903";
        when 902 => reg1_string <= " 902";
        when 901 => reg1_string <= " 901";
        when 900 => reg1_string <= " 900";
        when 899 => reg1_string <= " 899";
        when 898 => reg1_string <= " 898";
        when 897 => reg1_string <= " 897";
        when 896 => reg1_string <= " 896";
        when 895 => reg1_string <= " 895";
        when 894 => reg1_string <= " 894";
        when 893 => reg1_string <= " 893";
        when 892 => reg1_string <= " 892";
        when 891 => reg1_string <= " 891";
        when 890 => reg1_string <= " 890";
        when 889 => reg1_string <= " 889";
        when 888 => reg1_string <= " 888";
        when 887 => reg1_string <= " 887";
        when 886 => reg1_string <= " 886";
        when 885 => reg1_string <= " 885";
        when 884 => reg1_string <= " 884";
        when 883 => reg1_string <= " 883";
        when 882 => reg1_string <= " 882";
        when 881 => reg1_string <= " 881";
        when 880 => reg1_string <= " 880";
        when 879 => reg1_string <= " 879";
        when 878 => reg1_string <= " 878";
        when 877 => reg1_string <= " 877";
        when 876 => reg1_string <= " 876";
        when 875 => reg1_string <= " 875";
        when 874 => reg1_string <= " 874";
        when 873 => reg1_string <= " 873";
        when 872 => reg1_string <= " 872";
        when 871 => reg1_string <= " 871";
        when 870 => reg1_string <= " 870";
        when 869 => reg1_string <= " 869";
        when 868 => reg1_string <= " 868";
        when 867 => reg1_string <= " 867";
        when 866 => reg1_string <= " 866";
        when 865 => reg1_string <= " 865";
        when 864 => reg1_string <= " 864";
        when 863 => reg1_string <= " 863";
        when 862 => reg1_string <= " 862";
        when 861 => reg1_string <= " 861";
        when 860 => reg1_string <= " 860";
        when 859 => reg1_string <= " 859";
        when 858 => reg1_string <= " 858";
        when 857 => reg1_string <= " 857";
        when 856 => reg1_string <= " 856";
        when 855 => reg1_string <= " 855";
        when 854 => reg1_string <= " 854";
        when 853 => reg1_string <= " 853";
        when 852 => reg1_string <= " 852";
        when 851 => reg1_string <= " 851";
        when 850 => reg1_string <= " 850";
        when 849 => reg1_string <= " 849";
        when 848 => reg1_string <= " 848";
        when 847 => reg1_string <= " 847";
        when 846 => reg1_string <= " 846";
        when 845 => reg1_string <= " 845";
        when 844 => reg1_string <= " 844";
        when 843 => reg1_string <= " 843";
        when 842 => reg1_string <= " 842";
        when 841 => reg1_string <= " 841";
        when 840 => reg1_string <= " 840";
        when 839 => reg1_string <= " 839";
        when 838 => reg1_string <= " 838";
        when 837 => reg1_string <= " 837";
        when 836 => reg1_string <= " 836";
        when 835 => reg1_string <= " 835";
        when 834 => reg1_string <= " 834";
        when 833 => reg1_string <= " 833";
        when 832 => reg1_string <= " 832";
        when 831 => reg1_string <= " 831";
        when 830 => reg1_string <= " 830";
        when 829 => reg1_string <= " 829";
        when 828 => reg1_string <= " 828";
        when 827 => reg1_string <= " 827";
        when 826 => reg1_string <= " 826";
        when 825 => reg1_string <= " 825";
        when 824 => reg1_string <= " 824";
        when 823 => reg1_string <= " 823";
        when 822 => reg1_string <= " 822";
        when 821 => reg1_string <= " 821";
        when 820 => reg1_string <= " 820";
        when 819 => reg1_string <= " 819";
        when 818 => reg1_string <= " 818";
        when 817 => reg1_string <= " 817";
        when 816 => reg1_string <= " 816";
        when 815 => reg1_string <= " 815";
        when 814 => reg1_string <= " 814";
        when 813 => reg1_string <= " 813";
        when 812 => reg1_string <= " 812";
        when 811 => reg1_string <= " 811";
        when 810 => reg1_string <= " 810";
        when 809 => reg1_string <= " 809";
        when 808 => reg1_string <= " 808";
        when 807 => reg1_string <= " 807";
        when 806 => reg1_string <= " 806";
        when 805 => reg1_string <= " 805";
        when 804 => reg1_string <= " 804";
        when 803 => reg1_string <= " 803";
        when 802 => reg1_string <= " 802";
        when 801 => reg1_string <= " 801";
        when 800 => reg1_string <= " 800";
        when 799 => reg1_string <= " 799";
        when 798 => reg1_string <= " 798";
        when 797 => reg1_string <= " 797";
        when 796 => reg1_string <= " 796";
        when 795 => reg1_string <= " 795";
        when 794 => reg1_string <= " 794";
        when 793 => reg1_string <= " 793";
        when 792 => reg1_string <= " 792";
        when 791 => reg1_string <= " 791";
        when 790 => reg1_string <= " 790";
        when 789 => reg1_string <= " 789";
        when 788 => reg1_string <= " 788";
        when 787 => reg1_string <= " 787";
        when 786 => reg1_string <= " 786";
        when 785 => reg1_string <= " 785";
        when 784 => reg1_string <= " 784";
        when 783 => reg1_string <= " 783";
        when 782 => reg1_string <= " 782";
        when 781 => reg1_string <= " 781";
        when 780 => reg1_string <= " 780";
        when 779 => reg1_string <= " 779";
        when 778 => reg1_string <= " 778";
        when 777 => reg1_string <= " 777";
        when 776 => reg1_string <= " 776";
        when 775 => reg1_string <= " 775";
        when 774 => reg1_string <= " 774";
        when 773 => reg1_string <= " 773";
        when 772 => reg1_string <= " 772";
        when 771 => reg1_string <= " 771";
        when 770 => reg1_string <= " 770";
        when 769 => reg1_string <= " 769";
        when 768 => reg1_string <= " 768";
        when 767 => reg1_string <= " 767";
        when 766 => reg1_string <= " 766";
        when 765 => reg1_string <= " 765";
        when 764 => reg1_string <= " 764";
        when 763 => reg1_string <= " 763";
        when 762 => reg1_string <= " 762";
        when 761 => reg1_string <= " 761";
        when 760 => reg1_string <= " 760";
        when 759 => reg1_string <= " 759";
        when 758 => reg1_string <= " 758";
        when 757 => reg1_string <= " 757";
        when 756 => reg1_string <= " 756";
        when 755 => reg1_string <= " 755";
        when 754 => reg1_string <= " 754";
        when 753 => reg1_string <= " 753";
        when 752 => reg1_string <= " 752";
        when 751 => reg1_string <= " 751";
        when 750 => reg1_string <= " 750";
        when 749 => reg1_string <= " 749";
        when 748 => reg1_string <= " 748";
        when 747 => reg1_string <= " 747";
        when 746 => reg1_string <= " 746";
        when 745 => reg1_string <= " 745";
        when 744 => reg1_string <= " 744";
        when 743 => reg1_string <= " 743";
        when 742 => reg1_string <= " 742";
        when 741 => reg1_string <= " 741";
        when 740 => reg1_string <= " 740";
        when 739 => reg1_string <= " 739";
        when 738 => reg1_string <= " 738";
        when 737 => reg1_string <= " 737";
        when 736 => reg1_string <= " 736";
        when 735 => reg1_string <= " 735";
        when 734 => reg1_string <= " 734";
        when 733 => reg1_string <= " 733";
        when 732 => reg1_string <= " 732";
        when 731 => reg1_string <= " 731";
        when 730 => reg1_string <= " 730";
        when 729 => reg1_string <= " 729";
        when 728 => reg1_string <= " 728";
        when 727 => reg1_string <= " 727";
        when 726 => reg1_string <= " 726";
        when 725 => reg1_string <= " 725";
        when 724 => reg1_string <= " 724";
        when 723 => reg1_string <= " 723";
        when 722 => reg1_string <= " 722";
        when 721 => reg1_string <= " 721";
        when 720 => reg1_string <= " 720";
        when 719 => reg1_string <= " 719";
        when 718 => reg1_string <= " 718";
        when 717 => reg1_string <= " 717";
        when 716 => reg1_string <= " 716";
        when 715 => reg1_string <= " 715";
        when 714 => reg1_string <= " 714";
        when 713 => reg1_string <= " 713";
        when 712 => reg1_string <= " 712";
        when 711 => reg1_string <= " 711";
        when 710 => reg1_string <= " 710";
        when 709 => reg1_string <= " 709";
        when 708 => reg1_string <= " 708";
        when 707 => reg1_string <= " 707";
        when 706 => reg1_string <= " 706";
        when 705 => reg1_string <= " 705";
        when 704 => reg1_string <= " 704";
        when 703 => reg1_string <= " 703";
        when 702 => reg1_string <= " 702";
        when 701 => reg1_string <= " 701";
        when 700 => reg1_string <= " 700";
        when 699 => reg1_string <= " 699";
        when 698 => reg1_string <= " 698";
        when 697 => reg1_string <= " 697";
        when 696 => reg1_string <= " 696";
        when 695 => reg1_string <= " 695";
        when 694 => reg1_string <= " 694";
        when 693 => reg1_string <= " 693";
        when 692 => reg1_string <= " 692";
        when 691 => reg1_string <= " 691";
        when 690 => reg1_string <= " 690";
        when 689 => reg1_string <= " 689";
        when 688 => reg1_string <= " 688";
        when 687 => reg1_string <= " 687";
        when 686 => reg1_string <= " 686";
        when 685 => reg1_string <= " 685";
        when 684 => reg1_string <= " 684";
        when 683 => reg1_string <= " 683";
        when 682 => reg1_string <= " 682";
        when 681 => reg1_string <= " 681";
        when 680 => reg1_string <= " 680";
        when 679 => reg1_string <= " 679";
        when 678 => reg1_string <= " 678";
        when 677 => reg1_string <= " 677";
        when 676 => reg1_string <= " 676";
        when 675 => reg1_string <= " 675";
        when 674 => reg1_string <= " 674";
        when 673 => reg1_string <= " 673";
        when 672 => reg1_string <= " 672";
        when 671 => reg1_string <= " 671";
        when 670 => reg1_string <= " 670";
        when 669 => reg1_string <= " 669";
        when 668 => reg1_string <= " 668";
        when 667 => reg1_string <= " 667";
        when 666 => reg1_string <= " 666";
        when 665 => reg1_string <= " 665";
        when 664 => reg1_string <= " 664";
        when 663 => reg1_string <= " 663";
        when 662 => reg1_string <= " 662";
        when 661 => reg1_string <= " 661";
        when 660 => reg1_string <= " 660";
        when 659 => reg1_string <= " 659";
        when 658 => reg1_string <= " 658";
        when 657 => reg1_string <= " 657";
        when 656 => reg1_string <= " 656";
        when 655 => reg1_string <= " 655";
        when 654 => reg1_string <= " 654";
        when 653 => reg1_string <= " 653";
        when 652 => reg1_string <= " 652";
        when 651 => reg1_string <= " 651";
        when 650 => reg1_string <= " 650";
        when 649 => reg1_string <= " 649";
        when 648 => reg1_string <= " 648";
        when 647 => reg1_string <= " 647";
        when 646 => reg1_string <= " 646";
        when 645 => reg1_string <= " 645";
        when 644 => reg1_string <= " 644";
        when 643 => reg1_string <= " 643";
        when 642 => reg1_string <= " 642";
        when 641 => reg1_string <= " 641";
        when 640 => reg1_string <= " 640";
        when 639 => reg1_string <= " 639";
        when 638 => reg1_string <= " 638";
        when 637 => reg1_string <= " 637";
        when 636 => reg1_string <= " 636";
        when 635 => reg1_string <= " 635";
        when 634 => reg1_string <= " 634";
        when 633 => reg1_string <= " 633";
        when 632 => reg1_string <= " 632";
        when 631 => reg1_string <= " 631";
        when 630 => reg1_string <= " 630";
        when 629 => reg1_string <= " 629";
        when 628 => reg1_string <= " 628";
        when 627 => reg1_string <= " 627";
        when 626 => reg1_string <= " 626";
        when 625 => reg1_string <= " 625";
        when 624 => reg1_string <= " 624";
        when 623 => reg1_string <= " 623";
        when 622 => reg1_string <= " 622";
        when 621 => reg1_string <= " 621";
        when 620 => reg1_string <= " 620";
        when 619 => reg1_string <= " 619";
        when 618 => reg1_string <= " 618";
        when 617 => reg1_string <= " 617";
        when 616 => reg1_string <= " 616";
        when 615 => reg1_string <= " 615";
        when 614 => reg1_string <= " 614";
        when 613 => reg1_string <= " 613";
        when 612 => reg1_string <= " 612";
        when 611 => reg1_string <= " 611";
        when 610 => reg1_string <= " 610";
        when 609 => reg1_string <= " 609";
        when 608 => reg1_string <= " 608";
        when 607 => reg1_string <= " 607";
        when 606 => reg1_string <= " 606";
        when 605 => reg1_string <= " 605";
        when 604 => reg1_string <= " 604";
        when 603 => reg1_string <= " 603";
        when 602 => reg1_string <= " 602";
        when 601 => reg1_string <= " 601";
        when 600 => reg1_string <= " 600";
        when 599 => reg1_string <= " 599";
        when 598 => reg1_string <= " 598";
        when 597 => reg1_string <= " 597";
        when 596 => reg1_string <= " 596";
        when 595 => reg1_string <= " 595";
        when 594 => reg1_string <= " 594";
        when 593 => reg1_string <= " 593";
        when 592 => reg1_string <= " 592";
        when 591 => reg1_string <= " 591";
        when 590 => reg1_string <= " 590";
        when 589 => reg1_string <= " 589";
        when 588 => reg1_string <= " 588";
        when 587 => reg1_string <= " 587";
        when 586 => reg1_string <= " 586";
        when 585 => reg1_string <= " 585";
        when 584 => reg1_string <= " 584";
        when 583 => reg1_string <= " 583";
        when 582 => reg1_string <= " 582";
        when 581 => reg1_string <= " 581";
        when 580 => reg1_string <= " 580";
        when 579 => reg1_string <= " 579";
        when 578 => reg1_string <= " 578";
        when 577 => reg1_string <= " 577";
        when 576 => reg1_string <= " 576";
        when 575 => reg1_string <= " 575";
        when 574 => reg1_string <= " 574";
        when 573 => reg1_string <= " 573";
        when 572 => reg1_string <= " 572";
        when 571 => reg1_string <= " 571";
        when 570 => reg1_string <= " 570";
        when 569 => reg1_string <= " 569";
        when 568 => reg1_string <= " 568";
        when 567 => reg1_string <= " 567";
        when 566 => reg1_string <= " 566";
        when 565 => reg1_string <= " 565";
        when 564 => reg1_string <= " 564";
        when 563 => reg1_string <= " 563";
        when 562 => reg1_string <= " 562";
        when 561 => reg1_string <= " 561";
        when 560 => reg1_string <= " 560";
        when 559 => reg1_string <= " 559";
        when 558 => reg1_string <= " 558";
        when 557 => reg1_string <= " 557";
        when 556 => reg1_string <= " 556";
        when 555 => reg1_string <= " 555";
        when 554 => reg1_string <= " 554";
        when 553 => reg1_string <= " 553";
        when 552 => reg1_string <= " 552";
        when 551 => reg1_string <= " 551";
        when 550 => reg1_string <= " 550";
        when 549 => reg1_string <= " 549";
        when 548 => reg1_string <= " 548";
        when 547 => reg1_string <= " 547";
        when 546 => reg1_string <= " 546";
        when 545 => reg1_string <= " 545";
        when 544 => reg1_string <= " 544";
        when 543 => reg1_string <= " 543";
        when 542 => reg1_string <= " 542";
        when 541 => reg1_string <= " 541";
        when 540 => reg1_string <= " 540";
        when 539 => reg1_string <= " 539";
        when 538 => reg1_string <= " 538";
        when 537 => reg1_string <= " 537";
        when 536 => reg1_string <= " 536";
        when 535 => reg1_string <= " 535";
        when 534 => reg1_string <= " 534";
        when 533 => reg1_string <= " 533";
        when 532 => reg1_string <= " 532";
        when 531 => reg1_string <= " 531";
        when 530 => reg1_string <= " 530";
        when 529 => reg1_string <= " 529";
        when 528 => reg1_string <= " 528";
        when 527 => reg1_string <= " 527";
        when 526 => reg1_string <= " 526";
        when 525 => reg1_string <= " 525";
        when 524 => reg1_string <= " 524";
        when 523 => reg1_string <= " 523";
        when 522 => reg1_string <= " 522";
        when 521 => reg1_string <= " 521";
        when 520 => reg1_string <= " 520";
        when 519 => reg1_string <= " 519";
        when 518 => reg1_string <= " 518";
        when 517 => reg1_string <= " 517";
        when 516 => reg1_string <= " 516";
        when 515 => reg1_string <= " 515";
        when 514 => reg1_string <= " 514";
        when 513 => reg1_string <= " 513";
        when 512 => reg1_string <= " 512";
        when 511 => reg1_string <= " 511";
        when 510 => reg1_string <= " 510";
        when 509 => reg1_string <= " 509";
        when 508 => reg1_string <= " 508";
        when 507 => reg1_string <= " 507";
        when 506 => reg1_string <= " 506";
        when 505 => reg1_string <= " 505";
        when 504 => reg1_string <= " 504";
        when 503 => reg1_string <= " 503";
        when 502 => reg1_string <= " 502";
        when 501 => reg1_string <= " 501";
        when 500 => reg1_string <= " 500";
        when 499 => reg1_string <= " 499";
        when 498 => reg1_string <= " 498";
        when 497 => reg1_string <= " 497";
        when 496 => reg1_string <= " 496";
        when 495 => reg1_string <= " 495";
        when 494 => reg1_string <= " 494";
        when 493 => reg1_string <= " 493";
        when 492 => reg1_string <= " 492";
        when 491 => reg1_string <= " 491";
        when 490 => reg1_string <= " 490";
        when 489 => reg1_string <= " 489";
        when 488 => reg1_string <= " 488";
        when 487 => reg1_string <= " 487";
        when 486 => reg1_string <= " 486";
        when 485 => reg1_string <= " 485";
        when 484 => reg1_string <= " 484";
        when 483 => reg1_string <= " 483";
        when 482 => reg1_string <= " 482";
        when 481 => reg1_string <= " 481";
        when 480 => reg1_string <= " 480";
        when 479 => reg1_string <= " 479";
        when 478 => reg1_string <= " 478";
        when 477 => reg1_string <= " 477";
        when 476 => reg1_string <= " 476";
        when 475 => reg1_string <= " 475";
        when 474 => reg1_string <= " 474";
        when 473 => reg1_string <= " 473";
        when 472 => reg1_string <= " 472";
        when 471 => reg1_string <= " 471";
        when 470 => reg1_string <= " 470";
        when 469 => reg1_string <= " 469";
        when 468 => reg1_string <= " 468";
        when 467 => reg1_string <= " 467";
        when 466 => reg1_string <= " 466";
        when 465 => reg1_string <= " 465";
        when 464 => reg1_string <= " 464";
        when 463 => reg1_string <= " 463";
        when 462 => reg1_string <= " 462";
        when 461 => reg1_string <= " 461";
        when 460 => reg1_string <= " 460";
        when 459 => reg1_string <= " 459";
        when 458 => reg1_string <= " 458";
        when 457 => reg1_string <= " 457";
        when 456 => reg1_string <= " 456";
        when 455 => reg1_string <= " 455";
        when 454 => reg1_string <= " 454";
        when 453 => reg1_string <= " 453";
        when 452 => reg1_string <= " 452";
        when 451 => reg1_string <= " 451";
        when 450 => reg1_string <= " 450";
        when 449 => reg1_string <= " 449";
        when 448 => reg1_string <= " 448";
        when 447 => reg1_string <= " 447";
        when 446 => reg1_string <= " 446";
        when 445 => reg1_string <= " 445";
        when 444 => reg1_string <= " 444";
        when 443 => reg1_string <= " 443";
        when 442 => reg1_string <= " 442";
        when 441 => reg1_string <= " 441";
        when 440 => reg1_string <= " 440";
        when 439 => reg1_string <= " 439";
        when 438 => reg1_string <= " 438";
        when 437 => reg1_string <= " 437";
        when 436 => reg1_string <= " 436";
        when 435 => reg1_string <= " 435";
        when 434 => reg1_string <= " 434";
        when 433 => reg1_string <= " 433";
        when 432 => reg1_string <= " 432";
        when 431 => reg1_string <= " 431";
        when 430 => reg1_string <= " 430";
        when 429 => reg1_string <= " 429";
        when 428 => reg1_string <= " 428";
        when 427 => reg1_string <= " 427";
        when 426 => reg1_string <= " 426";
        when 425 => reg1_string <= " 425";
        when 424 => reg1_string <= " 424";
        when 423 => reg1_string <= " 423";
        when 422 => reg1_string <= " 422";
        when 421 => reg1_string <= " 421";
        when 420 => reg1_string <= " 420";
        when 419 => reg1_string <= " 419";
        when 418 => reg1_string <= " 418";
        when 417 => reg1_string <= " 417";
        when 416 => reg1_string <= " 416";
        when 415 => reg1_string <= " 415";
        when 414 => reg1_string <= " 414";
        when 413 => reg1_string <= " 413";
        when 412 => reg1_string <= " 412";
        when 411 => reg1_string <= " 411";
        when 410 => reg1_string <= " 410";
        when 409 => reg1_string <= " 409";
        when 408 => reg1_string <= " 408";
        when 407 => reg1_string <= " 407";
        when 406 => reg1_string <= " 406";
        when 405 => reg1_string <= " 405";
        when 404 => reg1_string <= " 404";
        when 403 => reg1_string <= " 403";
        when 402 => reg1_string <= " 402";
        when 401 => reg1_string <= " 401";
        when 400 => reg1_string <= " 400";
        when 399 => reg1_string <= " 399";
        when 398 => reg1_string <= " 398";
        when 397 => reg1_string <= " 397";
        when 396 => reg1_string <= " 396";
        when 395 => reg1_string <= " 395";
        when 394 => reg1_string <= " 394";
        when 393 => reg1_string <= " 393";
        when 392 => reg1_string <= " 392";
        when 391 => reg1_string <= " 391";
        when 390 => reg1_string <= " 390";
        when 389 => reg1_string <= " 389";
        when 388 => reg1_string <= " 388";
        when 387 => reg1_string <= " 387";
        when 386 => reg1_string <= " 386";
        when 385 => reg1_string <= " 385";
        when 384 => reg1_string <= " 384";
        when 383 => reg1_string <= " 383";
        when 382 => reg1_string <= " 382";
        when 381 => reg1_string <= " 381";
        when 380 => reg1_string <= " 380";
        when 379 => reg1_string <= " 379";
        when 378 => reg1_string <= " 378";
        when 377 => reg1_string <= " 377";
        when 376 => reg1_string <= " 376";
        when 375 => reg1_string <= " 375";
        when 374 => reg1_string <= " 374";
        when 373 => reg1_string <= " 373";
        when 372 => reg1_string <= " 372";
        when 371 => reg1_string <= " 371";
        when 370 => reg1_string <= " 370";
        when 369 => reg1_string <= " 369";
        when 368 => reg1_string <= " 368";
        when 367 => reg1_string <= " 367";
        when 366 => reg1_string <= " 366";
        when 365 => reg1_string <= " 365";
        when 364 => reg1_string <= " 364";
        when 363 => reg1_string <= " 363";
        when 362 => reg1_string <= " 362";
        when 361 => reg1_string <= " 361";
        when 360 => reg1_string <= " 360";
        when 359 => reg1_string <= " 359";
        when 358 => reg1_string <= " 358";
        when 357 => reg1_string <= " 357";
        when 356 => reg1_string <= " 356";
        when 355 => reg1_string <= " 355";
        when 354 => reg1_string <= " 354";
        when 353 => reg1_string <= " 353";
        when 352 => reg1_string <= " 352";
        when 351 => reg1_string <= " 351";
        when 350 => reg1_string <= " 350";
        when 349 => reg1_string <= " 349";
        when 348 => reg1_string <= " 348";
        when 347 => reg1_string <= " 347";
        when 346 => reg1_string <= " 346";
        when 345 => reg1_string <= " 345";
        when 344 => reg1_string <= " 344";
        when 343 => reg1_string <= " 343";
        when 342 => reg1_string <= " 342";
        when 341 => reg1_string <= " 341";
        when 340 => reg1_string <= " 340";
        when 339 => reg1_string <= " 339";
        when 338 => reg1_string <= " 338";
        when 337 => reg1_string <= " 337";
        when 336 => reg1_string <= " 336";
        when 335 => reg1_string <= " 335";
        when 334 => reg1_string <= " 334";
        when 333 => reg1_string <= " 333";
        when 332 => reg1_string <= " 332";
        when 331 => reg1_string <= " 331";
        when 330 => reg1_string <= " 330";
        when 329 => reg1_string <= " 329";
        when 328 => reg1_string <= " 328";
        when 327 => reg1_string <= " 327";
        when 326 => reg1_string <= " 326";
        when 325 => reg1_string <= " 325";
        when 324 => reg1_string <= " 324";
        when 323 => reg1_string <= " 323";
        when 322 => reg1_string <= " 322";
        when 321 => reg1_string <= " 321";
        when 320 => reg1_string <= " 320";
        when 319 => reg1_string <= " 319";
        when 318 => reg1_string <= " 318";
        when 317 => reg1_string <= " 317";
        when 316 => reg1_string <= " 316";
        when 315 => reg1_string <= " 315";
        when 314 => reg1_string <= " 314";
        when 313 => reg1_string <= " 313";
        when 312 => reg1_string <= " 312";
        when 311 => reg1_string <= " 311";
        when 310 => reg1_string <= " 310";
        when 309 => reg1_string <= " 309";
        when 308 => reg1_string <= " 308";
        when 307 => reg1_string <= " 307";
        when 306 => reg1_string <= " 306";
        when 305 => reg1_string <= " 305";
        when 304 => reg1_string <= " 304";
        when 303 => reg1_string <= " 303";
        when 302 => reg1_string <= " 302";
        when 301 => reg1_string <= " 301";
        when 300 => reg1_string <= " 300";
        when 299 => reg1_string <= " 299";
        when 298 => reg1_string <= " 298";
        when 297 => reg1_string <= " 297";
        when 296 => reg1_string <= " 296";
        when 295 => reg1_string <= " 295";
        when 294 => reg1_string <= " 294";
        when 293 => reg1_string <= " 293";
        when 292 => reg1_string <= " 292";
        when 291 => reg1_string <= " 291";
        when 290 => reg1_string <= " 290";
        when 289 => reg1_string <= " 289";
        when 288 => reg1_string <= " 288";
        when 287 => reg1_string <= " 287";
        when 286 => reg1_string <= " 286";
        when 285 => reg1_string <= " 285";
        when 284 => reg1_string <= " 284";
        when 283 => reg1_string <= " 283";
        when 282 => reg1_string <= " 282";
        when 281 => reg1_string <= " 281";
        when 280 => reg1_string <= " 280";
        when 279 => reg1_string <= " 279";
        when 278 => reg1_string <= " 278";
        when 277 => reg1_string <= " 277";
        when 276 => reg1_string <= " 276";
        when 275 => reg1_string <= " 275";
        when 274 => reg1_string <= " 274";
        when 273 => reg1_string <= " 273";
        when 272 => reg1_string <= " 272";
        when 271 => reg1_string <= " 271";
        when 270 => reg1_string <= " 270";
        when 269 => reg1_string <= " 269";
        when 268 => reg1_string <= " 268";
        when 267 => reg1_string <= " 267";
        when 266 => reg1_string <= " 266";
        when 265 => reg1_string <= " 265";
        when 264 => reg1_string <= " 264";
        when 263 => reg1_string <= " 263";
        when 262 => reg1_string <= " 262";
        when 261 => reg1_string <= " 261";
        when 260 => reg1_string <= " 260";
        when 259 => reg1_string <= " 259";
        when 258 => reg1_string <= " 258";
        when 257 => reg1_string <= " 257";
        when 256 => reg1_string <= " 256";
        when 255 => reg1_string <= " 255";
        when 254 => reg1_string <= " 254";
        when 253 => reg1_string <= " 253";
        when 252 => reg1_string <= " 252";
        when 251 => reg1_string <= " 251";
        when 250 => reg1_string <= " 250";
        when 249 => reg1_string <= " 249";
        when 248 => reg1_string <= " 248";
        when 247 => reg1_string <= " 247";
        when 246 => reg1_string <= " 246";
        when 245 => reg1_string <= " 245";
        when 244 => reg1_string <= " 244";
        when 243 => reg1_string <= " 243";
        when 242 => reg1_string <= " 242";
        when 241 => reg1_string <= " 241";
        when 240 => reg1_string <= " 240";
        when 239 => reg1_string <= " 239";
        when 238 => reg1_string <= " 238";
        when 237 => reg1_string <= " 237";
        when 236 => reg1_string <= " 236";
        when 235 => reg1_string <= " 235";
        when 234 => reg1_string <= " 234";
        when 233 => reg1_string <= " 233";
        when 232 => reg1_string <= " 232";
        when 231 => reg1_string <= " 231";
        when 230 => reg1_string <= " 230";
        when 229 => reg1_string <= " 229";
        when 228 => reg1_string <= " 228";
        when 227 => reg1_string <= " 227";
        when 226 => reg1_string <= " 226";
        when 225 => reg1_string <= " 225";
        when 224 => reg1_string <= " 224";
        when 223 => reg1_string <= " 223";
        when 222 => reg1_string <= " 222";
        when 221 => reg1_string <= " 221";
        when 220 => reg1_string <= " 220";
        when 219 => reg1_string <= " 219";
        when 218 => reg1_string <= " 218";
        when 217 => reg1_string <= " 217";
        when 216 => reg1_string <= " 216";
        when 215 => reg1_string <= " 215";
        when 214 => reg1_string <= " 214";
        when 213 => reg1_string <= " 213";
        when 212 => reg1_string <= " 212";
        when 211 => reg1_string <= " 211";
        when 210 => reg1_string <= " 210";
        when 209 => reg1_string <= " 209";
        when 208 => reg1_string <= " 208";
        when 207 => reg1_string <= " 207";
        when 206 => reg1_string <= " 206";
        when 205 => reg1_string <= " 205";
        when 204 => reg1_string <= " 204";
        when 203 => reg1_string <= " 203";
        when 202 => reg1_string <= " 202";
        when 201 => reg1_string <= " 201";
        when 200 => reg1_string <= " 200";
        when 199 => reg1_string <= " 199";
        when 198 => reg1_string <= " 198";
        when 197 => reg1_string <= " 197";
        when 196 => reg1_string <= " 196";
        when 195 => reg1_string <= " 195";
        when 194 => reg1_string <= " 194";
        when 193 => reg1_string <= " 193";
        when 192 => reg1_string <= " 192";
        when 191 => reg1_string <= " 191";
        when 190 => reg1_string <= " 190";
        when 189 => reg1_string <= " 189";
        when 188 => reg1_string <= " 188";
        when 187 => reg1_string <= " 187";
        when 186 => reg1_string <= " 186";
        when 185 => reg1_string <= " 185";
        when 184 => reg1_string <= " 184";
        when 183 => reg1_string <= " 183";
        when 182 => reg1_string <= " 182";
        when 181 => reg1_string <= " 181";
        when 180 => reg1_string <= " 180";
        when 179 => reg1_string <= " 179";
        when 178 => reg1_string <= " 178";
        when 177 => reg1_string <= " 177";
        when 176 => reg1_string <= " 176";
        when 175 => reg1_string <= " 175";
        when 174 => reg1_string <= " 174";
        when 173 => reg1_string <= " 173";
        when 172 => reg1_string <= " 172";
        when 171 => reg1_string <= " 171";
        when 170 => reg1_string <= " 170";
        when 169 => reg1_string <= " 169";
        when 168 => reg1_string <= " 168";
        when 167 => reg1_string <= " 167";
        when 166 => reg1_string <= " 166";
        when 165 => reg1_string <= " 165";
        when 164 => reg1_string <= " 164";
        when 163 => reg1_string <= " 163";
        when 162 => reg1_string <= " 162";
        when 161 => reg1_string <= " 161";
        when 160 => reg1_string <= " 160";
        when 159 => reg1_string <= " 159";
        when 158 => reg1_string <= " 158";
        when 157 => reg1_string <= " 157";
        when 156 => reg1_string <= " 156";
        when 155 => reg1_string <= " 155";
        when 154 => reg1_string <= " 154";
        when 153 => reg1_string <= " 153";
        when 152 => reg1_string <= " 152";
        when 151 => reg1_string <= " 151";
        when 150 => reg1_string <= " 150";
        when 149 => reg1_string <= " 149";
        when 148 => reg1_string <= " 148";
        when 147 => reg1_string <= " 147";
        when 146 => reg1_string <= " 146";
        when 145 => reg1_string <= " 145";
        when 144 => reg1_string <= " 144";
        when 143 => reg1_string <= " 143";
        when 142 => reg1_string <= " 142";
        when 141 => reg1_string <= " 141";
        when 140 => reg1_string <= " 140";
        when 139 => reg1_string <= " 139";
        when 138 => reg1_string <= " 138";
        when 137 => reg1_string <= " 137";
        when 136 => reg1_string <= " 136";
        when 135 => reg1_string <= " 135";
        when 134 => reg1_string <= " 134";
        when 133 => reg1_string <= " 133";
        when 132 => reg1_string <= " 132";
        when 131 => reg1_string <= " 131";
        when 130 => reg1_string <= " 130";
        when 129 => reg1_string <= " 129";
        when 128 => reg1_string <= " 128";
        when 127 => reg1_string <= " 127";
        when 126 => reg1_string <= " 126";
        when 125 => reg1_string <= " 125";
        when 124 => reg1_string <= " 124";
        when 123 => reg1_string <= " 123";
        when 122 => reg1_string <= " 122";
        when 121 => reg1_string <= " 121";
        when 120 => reg1_string <= " 120";
        when 119 => reg1_string <= " 119";
        when 118 => reg1_string <= " 118";
        when 117 => reg1_string <= " 117";
        when 116 => reg1_string <= " 116";
        when 115 => reg1_string <= " 115";
        when 114 => reg1_string <= " 114";
        when 113 => reg1_string <= " 113";
        when 112 => reg1_string <= " 112";
        when 111 => reg1_string <= " 111";
        when 110 => reg1_string <= " 110";
        when 109 => reg1_string <= " 109";
        when 108 => reg1_string <= " 108";
            when 107 => reg1_string <= " 107";                                                                                        
            when 106 => reg1_string <= " 106";                                                                                        
            when 105 => reg1_string <= " 105";                                                                                        
            when 104 => reg1_string <= " 104";                                                                                        
            when 103 => reg1_string <= " 103";                                                                                        
            when 102 => reg1_string <= " 102";                                                                                        
            when 101 => reg1_string <= " 101";                                                                                        
            when 100 => reg1_string <= " 100";                                                                                        
            when 99 => reg1_string <= "  99";                                                                                         
            when 98 => reg1_string <= "  98";                                                                                         
            when 97 => reg1_string <= "  97";                                                                                         
            when 96 => reg1_string <= "  96";                                                                                         
            when 95 => reg1_string <= "  95";                                                                                         
            when 94 => reg1_string <= "  94";                                                                                         
            when 93 => reg1_string <= "  93";                                                                                         
            when 92 => reg1_string <= "  92";                                                                                         
            when 91 => reg1_string <= "  91";                                                                                         
            when 90 => reg1_string <= "  90";                                                                                         
            when 89 => reg1_string <= "  89";                                                                                         
            when 88 => reg1_string <= "  88";                                                                                         
            when 87 => reg1_string <= "  87";                                                                                         
            when 86 => reg1_string <= "  86";                                                                                         
            when 85 => reg1_string <= "  85";                                                                                         
            when 84 => reg1_string <= "  84";                                                                                         
            when 83 => reg1_string <= "  83";                                                                                         
            when 82 => reg1_string <= "  82";                                                                                         
            when 81 => reg1_string <= "  81";                                                                                         
            when 80 => reg1_string <= "  80";                                                                                         
            when 79 => reg1_string <= "  79";                                                                                         
            when 78 => reg1_string <= "  78";                                                                                         
            when 77 => reg1_string <= "  77";
            when 76 => reg1_string <= "  76";                                                                                         
            when 75 => reg1_string <= "  75";                                                                                         
            when 74 => reg1_string <= "  74";                                                                                         
            when 73 => reg1_string <= "  73";                                                                                         
            when 72 => reg1_string <= "  72";                                                                                         
            when 71 => reg1_string <= "  71";                                                                                         
            when 70 => reg1_string <= "  70";                                                                                         
            when 69 => reg1_string <= "  69";                                                                                         
            when 68 => reg1_string <= "  68";                                                                                         
            when 67 => reg1_string <= "  67";                                                                                         
            when 66 => reg1_string <= "  66";                                                                                         
            when 65 => reg1_string <= "  65";                                                                                         
            when 64 => reg1_string <= "  64";                                                                                         
            when 63 => reg1_string <= "  63";                                                                                         
            when 62 => reg1_string <= "  62";                                                                                         
            when 61 => reg1_string <= "  61";                                                                                         
            when 60 => reg1_string <= "  60";                                                                                         
            when 59 => reg1_string <= "  59";                                                                                         
            when 58 => reg1_string <= "  58";                                                                                         
            when 57 => reg1_string <= "  57";                                                                                         
            when 56 => reg1_string <= "  56";                                                                                         
            when 55 => reg1_string <= "  55";                                                                                         
            when 54 => reg1_string <= "  54";                                                                                         
            when 53 => reg1_string <= "  53";                                                                                         
            when 52 => reg1_string <= "  52";                                                                                         
            when 51 => reg1_string <= "  51";                                                                                         
            when 50 => reg1_string <= "  50";                                                                                         
            when 49 => reg1_string <= "  49";                                                                                         
            when 48 => reg1_string <= "  48";                                                                                         
            when 47 => reg1_string <= "  47";
            when 46 => reg1_string <= "  46";                                                                                         
            when 45 => reg1_string <= "  45";                                                                                         
            when 44 => reg1_string <= "  44";                                                                                         
            when 43 => reg1_string <= "  43";                                                                                         
            when 42 => reg1_string <= "  42";                                                                                         
            when 41 => reg1_string <= "  41";                                                                                         
            when 40 => reg1_string <= "  40";                                                                                         
            when 39 => reg1_string <= "  39";                                                                                         
            when 38 => reg1_string <= "  38";                                                                                         
            when 37 => reg1_string <= "  37";                                                                                         
            when 36 => reg1_string <= "  36";                                                                                         
            when 35 => reg1_string <= "  35";                                                                                         
            when 34 => reg1_string <= "  34";                                                                                         
            when 33 => reg1_string <= "  33";                                                                                         
            when 32 => reg1_string <= "  32";                                                                                         
            when 31 => reg1_string <= "  31";                                                                                         
            when 30 => reg1_string <= "  30";                                                                                         
            when 29 => reg1_string <= "  29";                                                                                         
            when 28 => reg1_string <= "  28";                                                                                         
            when 27 => reg1_string <= "  27";                                                                                         
            when 26 => reg1_string <= "  26";                                                                                         
            when 25 => reg1_string <= "  25";                                                                                         
            when 24 => reg1_string <= "  24";                                                                                         
            when 23 => reg1_string <= "  23";
            when 22 => reg1_string <= "  22";                                                                                         
            when 21 => reg1_string <= "  21";                                                                                         
            when 20 => reg1_string <= "  20";                                                                                         
            when 19 => reg1_string <= "  19";                                                                                         
            when 18 => reg1_string <= "  18";                                                                                         
            when 17 => reg1_string <= "  17";                                                                                         
            when 16 => reg1_string <= "  16";                                                                                         
            when 15 => reg1_string <= "  15";                                                                                         
            when 14 => reg1_string <= "  14";                                                                                         
            when 13 => reg1_string <= "  13";                                                                                         
            when 12 => reg1_string <= "  12";                                                                                         
            when 11 => reg1_string <= "  11";                                                                                         
            when 10 => reg1_string <= "  10";                                                                                         
            when 9  => reg1_string <= "   9";                                                                                          
            when 8  => reg1_string <= "   8";                                                                                          
            when 7  => reg1_string <= "   7";                                                                                          
            when 6  => reg1_string <= "   6";                                                                                          
            when 5  => reg1_string <= "   5";                                                                                          
            when 4  => reg1_string <= "   4";                                                                                          
            when 3  => reg1_string <= "   3";                                                                                          
            when 2  => reg1_string <= "   2";                                                                                          
            when 1  => reg1_string <= "   1";                                                                                          
            when 0  => reg1_string <= "   0";
            when -1 => reg1_string <= "  -1";
            when -2 => reg1_string <= "  -2";
            when -3 => reg1_string <= "  -3";
            when -4 => reg1_string <= "  -4";
            when -5 => reg1_string <= "  -5";
            when -6 => reg1_string <= "  -6";
            when -7 => reg1_string <= "  -7";
            when -8 => reg1_string <= "  -8";
            when -9 => reg1_string <= "  -9";
            when -10 => reg1_string <= " -10";
            when -11 => reg1_string <= " -11";
            when -12 => reg1_string <= " -12";
            when -13 => reg1_string <= " -13";
            when -14 => reg1_string <= " -14";
            when -15 => reg1_string <= " -15";
            when -16 => reg1_string <= " -16";
            when -17 => reg1_string <= " -17";
            when -18 => reg1_string <= " -18";
            when -19 => reg1_string <= " -19";
            when -20 => reg1_string <= " -20";
            when -21 => reg1_string <= " -21";
            when -22 => reg1_string <= " -22";
            when -23 => reg1_string <= " -23";
            when -24 => reg1_string <= " -24";
            when -25 => reg1_string <= " -25";
            when -26 => reg1_string <= " -26";
            when -27 => reg1_string <= " -27";
            when -28 => reg1_string <= " -28";
            when -29 => reg1_string <= " -29";
            when -30 => reg1_string <= " -30";
            when -31 => reg1_string <= " -31";
            when -32 => reg1_string <= " -32";
            when -33 => reg1_string <= " -33";
            when -34 => reg1_string <= " -34";
            when -35 => reg1_string <= " -35";
            when -36 => reg1_string <= " -36";
            when -37 => reg1_string <= " -37";
            when -38 => reg1_string <= " -38";
            when -39 => reg1_string <= " -39";
            when -40 => reg1_string <= " -40";
            when -41 => reg1_string <= " -41";
            when -42 => reg1_string <= " -42";
            when -43 => reg1_string <= " -43";
            when -44 => reg1_string <= " -44";
            when -45 => reg1_string <= " -45";
            when -46 => reg1_string <= " -46";
            when -47 => reg1_string <= " -47";
            when -48 => reg1_string <= " -48";
            when -49 => reg1_string <= " -49";
            when -50 => reg1_string <= " -50";
            when -51 => reg1_string <= " -51";
            when -52 => reg1_string <= " -52";
            when -53 => reg1_string <= " -53";
            when -54 => reg1_string <= " -54";
            when -55 => reg1_string <= " -55";
            when -56 => reg1_string <= " -56";
            when -57 => reg1_string <= " -57";
            when -58 => reg1_string <= " -58";
            when -59 => reg1_string <= " -59";
            when -60 => reg1_string <= " -60";
            when -61 => reg1_string <= " -61";
            when -62 => reg1_string <= " -62";
            when -63 => reg1_string <= " -63";
            when -64 => reg1_string <= " -64";
            when -65 => reg1_string <= " -65";
            when -66 => reg1_string <= " -66";
            when -67 => reg1_string <= " -67";
            when -68 => reg1_string <= " -68";
            when -69 => reg1_string <= " -69";
            when -70 => reg1_string <= " -70";
            when -71 => reg1_string <= " -71";
            when -72 => reg1_string <= " -72";
            when -73 => reg1_string <= " -73";
            when -74 => reg1_string <= " -74";
            when -75 => reg1_string <= " -75";
            when -76 => reg1_string <= " -76";
            when -77 => reg1_string <= " -77";
            when -78 => reg1_string <= " -78";
            when -79 => reg1_string <= " -79";
            when -80 => reg1_string <= " -80";
            when -81 => reg1_string <= " -81";
            when -82 => reg1_string <= " -82";
            when -83 => reg1_string <= " -83";
            when -84 => reg1_string <= " -84";
            when -85 => reg1_string <= " -85";
            when -86 => reg1_string <= " -86";
            when -87 => reg1_string <= " -87";
            when -88 => reg1_string <= " -88";
            when -89 => reg1_string <= " -89";
            when -90 => reg1_string <= " -90";
            when -91 => reg1_string <= " -91";
            when -92 => reg1_string <= " -92";
            when -93 => reg1_string <= " -93";
            when -94 => reg1_string <= " -94";
            when -95 => reg1_string <= " -95";
            when -96 => reg1_string <= " -96";
            when -97 => reg1_string <= " -97";
            when -98 => reg1_string <= " -98";
            when -99 => reg1_string <= " -99";
            when -100 => reg1_string <= "-100";
            when -101 => reg1_string <= "-101";
            when -102 => reg1_string <= "-102";
            when -103 => reg1_string <= "-103";
            when -104 => reg1_string <= "-104";
            when -105 => reg1_string <= "-105";
            when -106 => reg1_string <= "-106";
            when -107 => reg1_string <= "-107";
            when -108 => reg1_string <= "-108";
            when -109 => reg1_string <= "-109";
            when -110 => reg1_string <= "-110";
            when -111 => reg1_string <= "-111";
            when -112 => reg1_string <= "-112";
            when -113 => reg1_string <= "-113";
            when -114 => reg1_string <= "-114";
            when -115 => reg1_string <= "-115";
            when -116 => reg1_string <= "-116";
            when -117 => reg1_string <= "-117";
            when -118 => reg1_string <= "-118";
            when -119 => reg1_string <= "-119";
            when -120 => reg1_string <= "-120";
            when -121 => reg1_string <= "-121";
            when -122 => reg1_string <= "-122";
            when -123 => reg1_string <= "-123";
            when -124 => reg1_string <= "-124";
            when -125 => reg1_string <= "-125";
            when -126 => reg1_string <= "-126";
            when -127 => reg1_string <= "-127";
            when -128 => reg1_string <= "-128";
            when -129 => reg1_string <= "-129";
            when -130 => reg1_string <= "-130";
            when -131 => reg1_string <= "-131";
            when -132 => reg1_string <= "-132";
            when -133 => reg1_string <= "-133";
            when -134 => reg1_string <= "-134";
            when -135 => reg1_string <= "-135";
            when -136 => reg1_string <= "-136";
            when -137 => reg1_string <= "-137";
            when -138 => reg1_string <= "-138";
            when -139 => reg1_string <= "-139";
            when -140 => reg1_string <= "-140";
            when -141 => reg1_string <= "-141";
            when -142 => reg1_string <= "-142";
            when -143 => reg1_string <= "-143";
            when -144 => reg1_string <= "-144";
            when -145 => reg1_string <= "-145";
            when -146 => reg1_string <= "-146";
            when -147 => reg1_string <= "-147";
            when -148 => reg1_string <= "-148";
            when -149 => reg1_string <= "-149";
            when -150 => reg1_string <= "-150";
            when -151 => reg1_string <= "-151";
            when -152 => reg1_string <= "-152";
            when -153 => reg1_string <= "-153";
            when -154 => reg1_string <= "-154";
            when -155 => reg1_string <= "-155";
            when -156 => reg1_string <= "-156";
            when -157 => reg1_string <= "-157";
            when -158 => reg1_string <= "-158";
            when -159 => reg1_string <= "-159";
            when -160 => reg1_string <= "-160";
            when -161 => reg1_string <= "-161";
            when -162 => reg1_string <= "-162";
            when -163 => reg1_string <= "-163";
            when -164 => reg1_string <= "-164";
            when -165 => reg1_string <= "-165";
            when -166 => reg1_string <= "-166";
            when -167 => reg1_string <= "-167";
            when -168 => reg1_string <= "-168";
            when -169 => reg1_string <= "-169";
            when -170 => reg1_string <= "-170";
            when -171 => reg1_string <= "-171";
            when -172 => reg1_string <= "-172";
            when -173 => reg1_string <= "-173";
            when -174 => reg1_string <= "-174";
            when -175 => reg1_string <= "-175";
            when -176 => reg1_string <= "-176";
            when -177 => reg1_string <= "-177";
            when -178 => reg1_string <= "-178";
            when -179 => reg1_string <= "-179";
            when -180 => reg1_string <= "-180";
            when -181 => reg1_string <= "-181";
            when -182 => reg1_string <= "-182";
            when -183 => reg1_string <= "-183";
            when -184 => reg1_string <= "-184";
            when -185 => reg1_string <= "-185";
            when -186 => reg1_string <= "-186";
            when -187 => reg1_string <= "-187";
            when -188 => reg1_string <= "-188";
            when -189 => reg1_string <= "-189";
            when -190 => reg1_string <= "-190";
            when -191 => reg1_string <= "-191";
            when -192 => reg1_string <= "-192";
            when -193 => reg1_string <= "-193";
            when -194 => reg1_string <= "-194";
            when -195 => reg1_string <= "-195";
            when -196 => reg1_string <= "-196";
            when -197 => reg1_string <= "-197";
            when -198 => reg1_string <= "-198";
            when -199 => reg1_string <= "-199";
            when -200 => reg1_string <= "-200";
            when -201 => reg1_string <= "-201";
            when -202 => reg1_string <= "-202";
            when -203 => reg1_string <= "-203";
            when -204 => reg1_string <= "-204";
            when -205 => reg1_string <= "-205";
            when -206 => reg1_string <= "-206";
            when -207 => reg1_string <= "-207";
            when -208 => reg1_string <= "-208";
            when -209 => reg1_string <= "-209";
            when -210 => reg1_string <= "-210";
            when -211 => reg1_string <= "-211";
            when -212 => reg1_string <= "-212";
            when -213 => reg1_string <= "-213";
            when -214 => reg1_string <= "-214";
            when -215 => reg1_string <= "-215";
            when -216 => reg1_string <= "-216";
            when -217 => reg1_string <= "-217";
            when -218 => reg1_string <= "-218";
            when -219 => reg1_string <= "-219";
            when -220 => reg1_string <= "-220";
            when -221 => reg1_string <= "-221";
            when -222 => reg1_string <= "-222";
            when -223 => reg1_string <= "-223";
            when -224 => reg1_string <= "-224";
            when -225 => reg1_string <= "-225";
            when -226 => reg1_string <= "-226";
            when -227 => reg1_string <= "-227";
            when -228 => reg1_string <= "-228";
            when -229 => reg1_string <= "-229";
            when -230 => reg1_string <= "-230";
            when -231 => reg1_string <= "-231";
            when -232 => reg1_string <= "-232";
            when -233 => reg1_string <= "-233";
            when -234 => reg1_string <= "-234";
            when -235 => reg1_string <= "-235";
            when -236 => reg1_string <= "-236";
            when -237 => reg1_string <= "-237";
            when -238 => reg1_string <= "-238";
            when -239 => reg1_string <= "-239";
            when -240 => reg1_string <= "-240";
            when -241 => reg1_string <= "-241";
            when -242 => reg1_string <= "-242";
            when -243 => reg1_string <= "-243";
            when -244 => reg1_string <= "-244";
            when -245 => reg1_string <= "-245";
            when -246 => reg1_string <= "-246";
            when -247 => reg1_string <= "-247";
            when -248 => reg1_string <= "-248";
            when -249 => reg1_string <= "-249";
            when -250 => reg1_string <= "-250";
            when -251 => reg1_string <= "-251";
            when -252 => reg1_string <= "-252";
            when -253 => reg1_string <= "-253";
            when -254 => reg1_string <= "-254";
            when -255 => reg1_string <= "-255";
            when -256 => reg1_string <= "-256";
            when -257 => reg1_string <= "-257";
            when -258 => reg1_string <= "-258";
            when -259 => reg1_string <= "-259";
            when -260 => reg1_string <= "-260";
            when -261 => reg1_string <= "-261";
            when -262 => reg1_string <= "-262";
            when -263 => reg1_string <= "-263";
            when -264 => reg1_string <= "-264";
            when -265 => reg1_string <= "-265";
            when -266 => reg1_string <= "-266";
            when -267 => reg1_string <= "-267";
            when -268 => reg1_string <= "-268";
            when -269 => reg1_string <= "-269";
            when -270 => reg1_string <= "-270";
            when -271 => reg1_string <= "-271";
            when -272 => reg1_string <= "-272";
            when -273 => reg1_string <= "-273";
            when -274 => reg1_string <= "-274";
            when -275 => reg1_string <= "-275";
            when -276 => reg1_string <= "-276";
            when -277 => reg1_string <= "-277";
            when -278 => reg1_string <= "-278";
            when -279 => reg1_string <= "-279";
            when -280 => reg1_string <= "-280";
            when -281 => reg1_string <= "-281";
            when -282 => reg1_string <= "-282";
            when -283 => reg1_string <= "-283";
            when -284 => reg1_string <= "-284";
            when -285 => reg1_string <= "-285";
            when -286 => reg1_string <= "-286";
            when -287 => reg1_string <= "-287";
            when -288 => reg1_string <= "-288";
            when -289 => reg1_string <= "-289";
            when -290 => reg1_string <= "-290";
            when -291 => reg1_string <= "-291";
            when -292 => reg1_string <= "-292";
            when -293 => reg1_string <= "-293";
            when -294 => reg1_string <= "-294";
            when -295 => reg1_string <= "-295";
            when -296 => reg1_string <= "-296";
            when -297 => reg1_string <= "-297";
            when -298 => reg1_string <= "-298";
            when -299 => reg1_string <= "-299";
            when -300 => reg1_string <= "-300";
            when -301 => reg1_string <= "-301";
            when -302 => reg1_string <= "-302";
            when -303 => reg1_string <= "-303";
            when -304 => reg1_string <= "-304";
            when -305 => reg1_string <= "-305";
            when -306 => reg1_string <= "-306";
            when -307 => reg1_string <= "-307";
            when -308 => reg1_string <= "-308";
            when -309 => reg1_string <= "-309";
            when -310 => reg1_string <= "-310";
            when -311 => reg1_string <= "-311";
            when -312 => reg1_string <= "-312";
            when -313 => reg1_string <= "-313";
            when -314 => reg1_string <= "-314";
            when -315 => reg1_string <= "-315";
            when -316 => reg1_string <= "-316";
            when -317 => reg1_string <= "-317";
            when -318 => reg1_string <= "-318";
            when -319 => reg1_string <= "-319";
            when -320 => reg1_string <= "-320";
            when -321 => reg1_string <= "-321";
            when -322 => reg1_string <= "-322";
            when -323 => reg1_string <= "-323";
            when -324 => reg1_string <= "-324";
            when -325 => reg1_string <= "-325";
            when -326 => reg1_string <= "-326";
            when -327 => reg1_string <= "-327";
            when -328 => reg1_string <= "-328";
            when -329 => reg1_string <= "-329";
            when -330 => reg1_string <= "-330";
            when -331 => reg1_string <= "-331";
            when -332 => reg1_string <= "-332";
            when -333 => reg1_string <= "-333";
            when -334 => reg1_string <= "-334";
            when -335 => reg1_string <= "-335";
            when -336 => reg1_string <= "-336";
            when -337 => reg1_string <= "-337";
            when -338 => reg1_string <= "-338";
            when -339 => reg1_string <= "-339";
            when -340 => reg1_string <= "-340";
            when -341 => reg1_string <= "-341";
            when -342 => reg1_string <= "-342";
            when -343 => reg1_string <= "-343";
            when -344 => reg1_string <= "-344";
            when -345 => reg1_string <= "-345";
            when -346 => reg1_string <= "-346";
            when -347 => reg1_string <= "-347";
            when -348 => reg1_string <= "-348";
            when -349 => reg1_string <= "-349";
            when -350 => reg1_string <= "-350";
            when -351 => reg1_string <= "-351";
            when -352 => reg1_string <= "-352";
            when -353 => reg1_string <= "-353";
            when -354 => reg1_string <= "-354";
            when -355 => reg1_string <= "-355";
            when -356 => reg1_string <= "-356";
            when -357 => reg1_string <= "-357";
            when -358 => reg1_string <= "-358";
            when -359 => reg1_string <= "-359";
            when -360 => reg1_string <= "-360";
            when -361 => reg1_string <= "-361";
            when -362 => reg1_string <= "-362";
            when -363 => reg1_string <= "-363";
            when -364 => reg1_string <= "-364";
            when -365 => reg1_string <= "-365";
            when -366 => reg1_string <= "-366";
            when -367 => reg1_string <= "-367";
            when -368 => reg1_string <= "-368";
            when -369 => reg1_string <= "-369";
            when -370 => reg1_string <= "-370";
            when -371 => reg1_string <= "-371";
            when -372 => reg1_string <= "-372";
            when -373 => reg1_string <= "-373";
            when -374 => reg1_string <= "-374";
            when -375 => reg1_string <= "-375";
            when -376 => reg1_string <= "-376";
            when -377 => reg1_string <= "-377";
            when -378 => reg1_string <= "-378";
            when -379 => reg1_string <= "-379";
            when -380 => reg1_string <= "-380";
            when -381 => reg1_string <= "-381";
            when -382 => reg1_string <= "-382";
            when -383 => reg1_string <= "-383";
            when -384 => reg1_string <= "-384";
            when -385 => reg1_string <= "-385";
            when -386 => reg1_string <= "-386";
            when -387 => reg1_string <= "-387";
            when -388 => reg1_string <= "-388";
            when -389 => reg1_string <= "-389";
            when -390 => reg1_string <= "-390";
            when -391 => reg1_string <= "-391";
            when -392 => reg1_string <= "-392";
            when -393 => reg1_string <= "-393";
            when -394 => reg1_string <= "-394";
            when -395 => reg1_string <= "-395";
            when -396 => reg1_string <= "-396";
            when -397 => reg1_string <= "-397";
            when -398 => reg1_string <= "-398";
            when -399 => reg1_string <= "-399";
            when -400 => reg1_string <= "-400";
            when -401 => reg1_string <= "-401";
            when -402 => reg1_string <= "-402";
            when -403 => reg1_string <= "-403";
            when -404 => reg1_string <= "-404";
            when -405 => reg1_string <= "-405";
            when -406 => reg1_string <= "-406";
            when -407 => reg1_string <= "-407";
            when -408 => reg1_string <= "-408";
            when -409 => reg1_string <= "-409";
            when -410 => reg1_string <= "-410";
            when -411 => reg1_string <= "-411";
            when -412 => reg1_string <= "-412";
            when -413 => reg1_string <= "-413";
            when -414 => reg1_string <= "-414";
            when -415 => reg1_string <= "-415";
            when -416 => reg1_string <= "-416";
            when -417 => reg1_string <= "-417";
            when -418 => reg1_string <= "-418";
            when -419 => reg1_string <= "-419";
            when -420 => reg1_string <= "-420";
            when -421 => reg1_string <= "-421";
            when -422 => reg1_string <= "-422";
            when -423 => reg1_string <= "-423";
            when -424 => reg1_string <= "-424";
            when -425 => reg1_string <= "-425";
            when -426 => reg1_string <= "-426";
            when -427 => reg1_string <= "-427";
            when -428 => reg1_string <= "-428";
            when -429 => reg1_string <= "-429";
            when -430 => reg1_string <= "-430";
            when -431 => reg1_string <= "-431";
            when -432 => reg1_string <= "-432";
            when -433 => reg1_string <= "-433";
            when -434 => reg1_string <= "-434";
            when -435 => reg1_string <= "-435";
            when -436 => reg1_string <= "-436";
            when -437 => reg1_string <= "-437";
            when -438 => reg1_string <= "-438";
            when -439 => reg1_string <= "-439";
            when -440 => reg1_string <= "-440";
            when -441 => reg1_string <= "-441";
            when -442 => reg1_string <= "-442";
            when -443 => reg1_string <= "-443";
            when -444 => reg1_string <= "-444";
            when -445 => reg1_string <= "-445";
            when -446 => reg1_string <= "-446";
            when -447 => reg1_string <= "-447";
            when -448 => reg1_string <= "-448";
            when -449 => reg1_string <= "-449";
            when -450 => reg1_string <= "-450";
            when -451 => reg1_string <= "-451";
            when -452 => reg1_string <= "-452";
            when -453 => reg1_string <= "-453";
            when -454 => reg1_string <= "-454";
            when -455 => reg1_string <= "-455";
            when -456 => reg1_string <= "-456";
            when -457 => reg1_string <= "-457";
            when -458 => reg1_string <= "-458";
            when -459 => reg1_string <= "-459";
            when -460 => reg1_string <= "-460";
            when -461 => reg1_string <= "-461";
            when -462 => reg1_string <= "-462";
            when -463 => reg1_string <= "-463";
            when -464 => reg1_string <= "-464";
            when -465 => reg1_string <= "-465";
            when -466 => reg1_string <= "-466";
            when -467 => reg1_string <= "-467";
            when -468 => reg1_string <= "-468";
            when -469 => reg1_string <= "-469";
            when -470 => reg1_string <= "-470";
            when -471 => reg1_string <= "-471";
            when -472 => reg1_string <= "-472";
            when -473 => reg1_string <= "-473";
            when -474 => reg1_string <= "-474";
            when -475 => reg1_string <= "-475";
            when -476 => reg1_string <= "-476";
            when -477 => reg1_string <= "-477";
            when -478 => reg1_string <= "-478";
            when -479 => reg1_string <= "-479";
            when -480 => reg1_string <= "-480";
            when -481 => reg1_string <= "-481";
            when -482 => reg1_string <= "-482";
            when -483 => reg1_string <= "-483";
            when -484 => reg1_string <= "-484";
            when -485 => reg1_string <= "-485";
            when -486 => reg1_string <= "-486";
            when -487 => reg1_string <= "-487";
            when -488 => reg1_string <= "-488";
            when -489 => reg1_string <= "-489";
            when -490 => reg1_string <= "-490";
            when -491 => reg1_string <= "-491";
            when -492 => reg1_string <= "-492";
            when -493 => reg1_string <= "-493";
            when -494 => reg1_string <= "-494";
            when -495 => reg1_string <= "-495";
            when -496 => reg1_string <= "-496";
            when -497 => reg1_string <= "-497";
            when -498 => reg1_string <= "-498";
            when -499 => reg1_string <= "-499";
            when -500 => reg1_string <= "-500";
            when -501 => reg1_string <= "-501";
            when -502 => reg1_string <= "-502";
            when -503 => reg1_string <= "-503";
            when -504 => reg1_string <= "-504";
            when -505 => reg1_string <= "-505";
            when -506 => reg1_string <= "-506";
            when -507 => reg1_string <= "-507";
            when -508 => reg1_string <= "-508";
            when -509 => reg1_string <= "-509";
            when -510 => reg1_string <= "-510";
            when -511 => reg1_string <= "-511";
            when -512 => reg1_string <= "-512";
            when -513 => reg1_string <= "-513";
            when -514 => reg1_string <= "-514";
            when -515 => reg1_string <= "-515";
            when -516 => reg1_string <= "-516";
            when -517 => reg1_string <= "-517";
            when -518 => reg1_string <= "-518";
            when -519 => reg1_string <= "-519";
            when -520 => reg1_string <= "-520";
            when -521 => reg1_string <= "-521";
            when -522 => reg1_string <= "-522";
            when -523 => reg1_string <= "-523";
            when -524 => reg1_string <= "-524";
            when -525 => reg1_string <= "-525";
            when -526 => reg1_string <= "-526";
            when -527 => reg1_string <= "-527";
            when -528 => reg1_string <= "-528";
            when -529 => reg1_string <= "-529";
            when -530 => reg1_string <= "-530";
            when -531 => reg1_string <= "-531";
            when -532 => reg1_string <= "-532";
            when -533 => reg1_string <= "-533";
            when -534 => reg1_string <= "-534";
            when -535 => reg1_string <= "-535";
            when -536 => reg1_string <= "-536";
            when -537 => reg1_string <= "-537";
            when -538 => reg1_string <= "-538";
            when -539 => reg1_string <= "-539";
            when -540 => reg1_string <= "-540";
            when -541 => reg1_string <= "-541";
            when -542 => reg1_string <= "-542";
            when -543 => reg1_string <= "-543";
            when -544 => reg1_string <= "-544";
            when -545 => reg1_string <= "-545";
            when -546 => reg1_string <= "-546";
            when -547 => reg1_string <= "-547";
            when -548 => reg1_string <= "-548";
            when -549 => reg1_string <= "-549";
            when -550 => reg1_string <= "-550";
            when -551 => reg1_string <= "-551";
            when -552 => reg1_string <= "-552";
            when -553 => reg1_string <= "-553";
            when -554 => reg1_string <= "-554";
            when -555 => reg1_string <= "-555";
            when -556 => reg1_string <= "-556";
            when -557 => reg1_string <= "-557";
            when -558 => reg1_string <= "-558";
            when -559 => reg1_string <= "-559";
            when -560 => reg1_string <= "-560";
            when -561 => reg1_string <= "-561";
            when -562 => reg1_string <= "-562";
            when -563 => reg1_string <= "-563";
            when -564 => reg1_string <= "-564";
            when -565 => reg1_string <= "-565";
            when -566 => reg1_string <= "-566";
            when -567 => reg1_string <= "-567";
            when -568 => reg1_string <= "-568";
            when -569 => reg1_string <= "-569";
            when -570 => reg1_string <= "-570";
            when -571 => reg1_string <= "-571";
            when -572 => reg1_string <= "-572";
            when -573 => reg1_string <= "-573";
            when -574 => reg1_string <= "-574";
            when -575 => reg1_string <= "-575";
            when -576 => reg1_string <= "-576";
            when -577 => reg1_string <= "-577";
            when -578 => reg1_string <= "-578";
            when -579 => reg1_string <= "-579";
            when -580 => reg1_string <= "-580";
            when -581 => reg1_string <= "-581";
            when -582 => reg1_string <= "-582";
            when -583 => reg1_string <= "-583";
            when -584 => reg1_string <= "-584";
            when -585 => reg1_string <= "-585";
            when -586 => reg1_string <= "-586";
            when -587 => reg1_string <= "-587";
            when -588 => reg1_string <= "-588";
            when -589 => reg1_string <= "-589";
            when -590 => reg1_string <= "-590";
            when -591 => reg1_string <= "-591";
            when -592 => reg1_string <= "-592";
            when -593 => reg1_string <= "-593";
            when -594 => reg1_string <= "-594";
            when -595 => reg1_string <= "-595";
            when -596 => reg1_string <= "-596";
            when -597 => reg1_string <= "-597";
            when -598 => reg1_string <= "-598";
            when -599 => reg1_string <= "-599";
            when -600 => reg1_string <= "-600";
            when -601 => reg1_string <= "-601";
            when -602 => reg1_string <= "-602";
            when -603 => reg1_string <= "-603";
            when -604 => reg1_string <= "-604";
            when -605 => reg1_string <= "-605";
            when -606 => reg1_string <= "-606";
            when -607 => reg1_string <= "-607";
            when -608 => reg1_string <= "-608";
            when -609 => reg1_string <= "-609";
            when -610 => reg1_string <= "-610";
            when -611 => reg1_string <= "-611";
            when -612 => reg1_string <= "-612";
            when -613 => reg1_string <= "-613";
            when -614 => reg1_string <= "-614";
            when -615 => reg1_string <= "-615";
            when -616 => reg1_string <= "-616";
            when -617 => reg1_string <= "-617";
            when -618 => reg1_string <= "-618";
            when -619 => reg1_string <= "-619";
            when -620 => reg1_string <= "-620";
            when -621 => reg1_string <= "-621";
            when -622 => reg1_string <= "-622";
            when -623 => reg1_string <= "-623";
            when -624 => reg1_string <= "-624";
            when -625 => reg1_string <= "-625";
            when -626 => reg1_string <= "-626";
            when -627 => reg1_string <= "-627";
            when -628 => reg1_string <= "-628";
            when -629 => reg1_string <= "-629";
            when -630 => reg1_string <= "-630";
            when -631 => reg1_string <= "-631";
            when -632 => reg1_string <= "-632";
            when -633 => reg1_string <= "-633";
            when -634 => reg1_string <= "-634";
            when -635 => reg1_string <= "-635";
            when -636 => reg1_string <= "-636";
            when -637 => reg1_string <= "-637";
            when -638 => reg1_string <= "-638";
            when -639 => reg1_string <= "-639";
            when -640 => reg1_string <= "-640";
            when -641 => reg1_string <= "-641";
            when -642 => reg1_string <= "-642";
            when -643 => reg1_string <= "-643";
            when -644 => reg1_string <= "-644";
            when -645 => reg1_string <= "-645";
            when -646 => reg1_string <= "-646";
            when -647 => reg1_string <= "-647";
            when -648 => reg1_string <= "-648";
            when -649 => reg1_string <= "-649";
            when -650 => reg1_string <= "-650";
            when -651 => reg1_string <= "-651";
            when -652 => reg1_string <= "-652";
            when -653 => reg1_string <= "-653";
            when -654 => reg1_string <= "-654";
            when -655 => reg1_string <= "-655";
            when -656 => reg1_string <= "-656";
            when -657 => reg1_string <= "-657";
            when -658 => reg1_string <= "-658";
            when -659 => reg1_string <= "-659";
            when -660 => reg1_string <= "-660";
            when -661 => reg1_string <= "-661";
            when -662 => reg1_string <= "-662";
            when -663 => reg1_string <= "-663";
            when -664 => reg1_string <= "-664";
            when -665 => reg1_string <= "-665";
            when -666 => reg1_string <= "-666";
            when -667 => reg1_string <= "-667";
            when -668 => reg1_string <= "-668";
            when -669 => reg1_string <= "-669";
            when -670 => reg1_string <= "-670";
            when -671 => reg1_string <= "-671";
            when -672 => reg1_string <= "-672";
            when -673 => reg1_string <= "-673";
            when -674 => reg1_string <= "-674";
            when -675 => reg1_string <= "-675";
            when -676 => reg1_string <= "-676";
            when -677 => reg1_string <= "-677";
            when -678 => reg1_string <= "-678";
            when -679 => reg1_string <= "-679";
            when -680 => reg1_string <= "-680";
            when -681 => reg1_string <= "-681";
            when -682 => reg1_string <= "-682";
            when -683 => reg1_string <= "-683";
            when -684 => reg1_string <= "-684";
            when -685 => reg1_string <= "-685";
            when -686 => reg1_string <= "-686";
            when -687 => reg1_string <= "-687";
            when -688 => reg1_string <= "-688";
            when -689 => reg1_string <= "-689";
            when -690 => reg1_string <= "-690";
            when -691 => reg1_string <= "-691";
            when -692 => reg1_string <= "-692";
            when -693 => reg1_string <= "-693";
            when -694 => reg1_string <= "-694";
            when -695 => reg1_string <= "-695";
            when -696 => reg1_string <= "-696";
            when -697 => reg1_string <= "-697";
            when -698 => reg1_string <= "-698";
            when -699 => reg1_string <= "-699";
            when -700 => reg1_string <= "-700";
            when -701 => reg1_string <= "-701";
            when -702 => reg1_string <= "-702";
            when -703 => reg1_string <= "-703";
            when -704 => reg1_string <= "-704";
            when -705 => reg1_string <= "-705";
            when -706 => reg1_string <= "-706";
            when -707 => reg1_string <= "-707";
            when -708 => reg1_string <= "-708";
            when -709 => reg1_string <= "-709";
            when -710 => reg1_string <= "-710";
            when -711 => reg1_string <= "-711";
            when -712 => reg1_string <= "-712";
            when -713 => reg1_string <= "-713";
            when -714 => reg1_string <= "-714";
            when -715 => reg1_string <= "-715";
            when -716 => reg1_string <= "-716";
            when -717 => reg1_string <= "-717";
            when -718 => reg1_string <= "-718";
            when -719 => reg1_string <= "-719";
            when -720 => reg1_string <= "-720";
            when -721 => reg1_string <= "-721";
            when -722 => reg1_string <= "-722";
            when -723 => reg1_string <= "-723";
            when -724 => reg1_string <= "-724";
            when -725 => reg1_string <= "-725";
            when -726 => reg1_string <= "-726";
            when -727 => reg1_string <= "-727";
            when -728 => reg1_string <= "-728";
            when -729 => reg1_string <= "-729";
            when -730 => reg1_string <= "-730";
            when -731 => reg1_string <= "-731";
            when -732 => reg1_string <= "-732";
            when -733 => reg1_string <= "-733";
            when -734 => reg1_string <= "-734";
            when -735 => reg1_string <= "-735";
            when -736 => reg1_string <= "-736";
            when -737 => reg1_string <= "-737";
            when -738 => reg1_string <= "-738";
            when -739 => reg1_string <= "-739";
            when -740 => reg1_string <= "-740";
            when -741 => reg1_string <= "-741";
            when -742 => reg1_string <= "-742";
            when -743 => reg1_string <= "-743";
            when -744 => reg1_string <= "-744";
            when -745 => reg1_string <= "-745";
            when -746 => reg1_string <= "-746";
            when -747 => reg1_string <= "-747";
            when -748 => reg1_string <= "-748";
            when -749 => reg1_string <= "-749";
            when -750 => reg1_string <= "-750";
            when -751 => reg1_string <= "-751";
            when -752 => reg1_string <= "-752";
            when -753 => reg1_string <= "-753";
            when -754 => reg1_string <= "-754";
            when -755 => reg1_string <= "-755";
            when -756 => reg1_string <= "-756";
            when -757 => reg1_string <= "-757";
            when -758 => reg1_string <= "-758";
            when -759 => reg1_string <= "-759";
            when -760 => reg1_string <= "-760";
            when -761 => reg1_string <= "-761";
            when -762 => reg1_string <= "-762";
            when -763 => reg1_string <= "-763";
            when -764 => reg1_string <= "-764";
            when -765 => reg1_string <= "-765";
            when -766 => reg1_string <= "-766";
            when -767 => reg1_string <= "-767";
            when -768 => reg1_string <= "-768";
            when -769 => reg1_string <= "-769";
            when -770 => reg1_string <= "-770";
            when -771 => reg1_string <= "-771";
            when -772 => reg1_string <= "-772";
            when -773 => reg1_string <= "-773";
            when -774 => reg1_string <= "-774";
            when -775 => reg1_string <= "-775";
            when -776 => reg1_string <= "-776";
            when -777 => reg1_string <= "-777";
            when -778 => reg1_string <= "-778";
            when -779 => reg1_string <= "-779";
            when -780 => reg1_string <= "-780";
            when -781 => reg1_string <= "-781";
            when -782 => reg1_string <= "-782";
            when -783 => reg1_string <= "-783";
            when -784 => reg1_string <= "-784";
            when -785 => reg1_string <= "-785";
            when -786 => reg1_string <= "-786";
            when -787 => reg1_string <= "-787";
            when -788 => reg1_string <= "-788";
            when -789 => reg1_string <= "-789";
            when -790 => reg1_string <= "-790";
            when -791 => reg1_string <= "-791";
            when -792 => reg1_string <= "-792";
            when -793 => reg1_string <= "-793";
            when -794 => reg1_string <= "-794";
            when -795 => reg1_string <= "-795";
            when -796 => reg1_string <= "-796";
            when -797 => reg1_string <= "-797";
            when -798 => reg1_string <= "-798";
            when -799 => reg1_string <= "-799";
            when -800 => reg1_string <= "-800";
            when -801 => reg1_string <= "-801";
            when -802 => reg1_string <= "-802";
            when -803 => reg1_string <= "-803";
            when -804 => reg1_string <= "-804";
            when -805 => reg1_string <= "-805";
            when -806 => reg1_string <= "-806";
            when -807 => reg1_string <= "-807";
            when -808 => reg1_string <= "-808";
            when -809 => reg1_string <= "-809";
            when -810 => reg1_string <= "-810";
            when -811 => reg1_string <= "-811";
            when -812 => reg1_string <= "-812";
            when -813 => reg1_string <= "-813";
            when -814 => reg1_string <= "-814";
            when -815 => reg1_string <= "-815";
            when -816 => reg1_string <= "-816";
            when -817 => reg1_string <= "-817";
            when -818 => reg1_string <= "-818";
            when -819 => reg1_string <= "-819";
            when -820 => reg1_string <= "-820";
            when -821 => reg1_string <= "-821";
            when -822 => reg1_string <= "-822";
            when -823 => reg1_string <= "-823";
            when -824 => reg1_string <= "-824";
            when -825 => reg1_string <= "-825";
            when -826 => reg1_string <= "-826";
            when -827 => reg1_string <= "-827";
            when -828 => reg1_string <= "-828";
            when -829 => reg1_string <= "-829";
            when -830 => reg1_string <= "-830";
            when -831 => reg1_string <= "-831";
            when -832 => reg1_string <= "-832";
            when -833 => reg1_string <= "-833";
            when -834 => reg1_string <= "-834";
            when -835 => reg1_string <= "-835";
            when -836 => reg1_string <= "-836";
            when -837 => reg1_string <= "-837";
            when -838 => reg1_string <= "-838";
            when -839 => reg1_string <= "-839";
            when -840 => reg1_string <= "-840";
            when -841 => reg1_string <= "-841";
            when -842 => reg1_string <= "-842";
            when -843 => reg1_string <= "-843";
            when -844 => reg1_string <= "-844";
            when -845 => reg1_string <= "-845";
            when -846 => reg1_string <= "-846";
            when -847 => reg1_string <= "-847";
            when -848 => reg1_string <= "-848";
            when -849 => reg1_string <= "-849";
            when -850 => reg1_string <= "-850";
            when -851 => reg1_string <= "-851";
            when -852 => reg1_string <= "-852";
            when -853 => reg1_string <= "-853";
            when -854 => reg1_string <= "-854";
            when -855 => reg1_string <= "-855";
            when -856 => reg1_string <= "-856";
            when -857 => reg1_string <= "-857";
            when -858 => reg1_string <= "-858";
            when -859 => reg1_string <= "-859";
            when -860 => reg1_string <= "-860";
            when -861 => reg1_string <= "-861";
            when -862 => reg1_string <= "-862";
            when -863 => reg1_string <= "-863";
            when -864 => reg1_string <= "-864";
            when -865 => reg1_string <= "-865";
            when -866 => reg1_string <= "-866";
            when -867 => reg1_string <= "-867";
            when -868 => reg1_string <= "-868";
            when -869 => reg1_string <= "-869";
            when -870 => reg1_string <= "-870";
            when -871 => reg1_string <= "-871";
            when -872 => reg1_string <= "-872";
            when -873 => reg1_string <= "-873";
            when -874 => reg1_string <= "-874";
            when -875 => reg1_string <= "-875";
            when -876 => reg1_string <= "-876";
            when -877 => reg1_string <= "-877";
            when -878 => reg1_string <= "-878";
            when -879 => reg1_string <= "-879";
            when -880 => reg1_string <= "-880";
            when -881 => reg1_string <= "-881";
            when -882 => reg1_string <= "-882";
            when -883 => reg1_string <= "-883";
            when -884 => reg1_string <= "-884";
            when -885 => reg1_string <= "-885";
            when -886 => reg1_string <= "-886";
            when -887 => reg1_string <= "-887";
            when -888 => reg1_string <= "-888";
            when -889 => reg1_string <= "-889";
            when -890 => reg1_string <= "-890";
            when -891 => reg1_string <= "-891";
            when -892 => reg1_string <= "-892";
            when -893 => reg1_string <= "-893";
            when -894 => reg1_string <= "-894";
            when -895 => reg1_string <= "-895";
            when -896 => reg1_string <= "-896";
            when -897 => reg1_string <= "-897";
            when -898 => reg1_string <= "-898";
            when -899 => reg1_string <= "-899";
            when -900 => reg1_string <= "-900";
            when -901 => reg1_string <= "-901";
            when -902 => reg1_string <= "-902";
            when -903 => reg1_string <= "-903";
            when -904 => reg1_string <= "-904";
            when -905 => reg1_string <= "-905";
            when -906 => reg1_string <= "-906";
            when -907 => reg1_string <= "-907";
            when -908 => reg1_string <= "-908";
            when -909 => reg1_string <= "-909";
            when -910 => reg1_string <= "-910";
            when -911 => reg1_string <= "-911";
            when -912 => reg1_string <= "-912";
            when -913 => reg1_string <= "-913";
            when -914 => reg1_string <= "-914";
            when -915 => reg1_string <= "-915";
            when -916 => reg1_string <= "-916";
            when -917 => reg1_string <= "-917";
            when -918 => reg1_string <= "-918";
            when -919 => reg1_string <= "-919";
            when -920 => reg1_string <= "-920";
            when -921 => reg1_string <= "-921";
            when -922 => reg1_string <= "-922";
            when -923 => reg1_string <= "-923";
            when -924 => reg1_string <= "-924";
            when -925 => reg1_string <= "-925";
            when -926 => reg1_string <= "-926";
            when -927 => reg1_string <= "-927";
            when -928 => reg1_string <= "-928";
            when -929 => reg1_string <= "-929";
            when -930 => reg1_string <= "-930";
            when -931 => reg1_string <= "-931";
            when -932 => reg1_string <= "-932";
            when -933 => reg1_string <= "-933";
            when -934 => reg1_string <= "-934";
            when -935 => reg1_string <= "-935";
            when -936 => reg1_string <= "-936";
            when -937 => reg1_string <= "-937";
            when -938 => reg1_string <= "-938";
            when -939 => reg1_string <= "-939";
            when -940 => reg1_string <= "-940";
            when -941 => reg1_string <= "-941";
            when -942 => reg1_string <= "-942";
            when -943 => reg1_string <= "-943";
            when -944 => reg1_string <= "-944";
            when -945 => reg1_string <= "-945";
            when -946 => reg1_string <= "-946";
            when -947 => reg1_string <= "-947";
            when -948 => reg1_string <= "-948";
            when -949 => reg1_string <= "-949";
            when -950 => reg1_string <= "-950";
            when -951 => reg1_string <= "-951";
            when -952 => reg1_string <= "-952";
            when -953 => reg1_string <= "-953";
            when -954 => reg1_string <= "-954";
            when -955 => reg1_string <= "-955";
            when -956 => reg1_string <= "-956";
            when -957 => reg1_string <= "-957";
            when -958 => reg1_string <= "-958";
            when -959 => reg1_string <= "-959";
            when -960 => reg1_string <= "-960";
            when -961 => reg1_string <= "-961";
            when -962 => reg1_string <= "-962";
            when -963 => reg1_string <= "-963";
            when -964 => reg1_string <= "-964";
            when -965 => reg1_string <= "-965";
            when -966 => reg1_string <= "-966";
            when -967 => reg1_string <= "-967";
            when -968 => reg1_string <= "-968";
            when -969 => reg1_string <= "-969";
            when -970 => reg1_string <= "-970";
            when -971 => reg1_string <= "-971";
            when -972 => reg1_string <= "-972";
            when -973 => reg1_string <= "-973";
            when -974 => reg1_string <= "-974";
            when -975 => reg1_string <= "-975";
            when -976 => reg1_string <= "-976";
            when -977 => reg1_string <= "-977";
            when -978 => reg1_string <= "-978";
            when -979 => reg1_string <= "-979";
            when -980 => reg1_string <= "-980";
            when -981 => reg1_string <= "-981";
            when -982 => reg1_string <= "-982";
            when -983 => reg1_string <= "-983";
            when -984 => reg1_string <= "-984";
            when -985 => reg1_string <= "-985";
            when -986 => reg1_string <= "-986";
            when -987 => reg1_string <= "-987";
            when -988 => reg1_string <= "-988";
            when -989 => reg1_string <= "-989";
            when -990 => reg1_string <= "-990";
            when -991 => reg1_string <= "-991";
            when -992 => reg1_string <= "-992";
            when -993 => reg1_string <= "-993";
            when -994 => reg1_string <= "-994";
            when -995 => reg1_string <= "-995";
            when -996 => reg1_string <= "-996";
            when -997 => reg1_string <= "-997";
            when -998 => reg1_string <= "-998";
            when -999 => reg1_string <= "-999";
            when others => reg1_string <= "    ";
        end case;
        
        case (reg0_int) is 
                when 999 => reg0_string <= " 999";
            when 998 => reg0_string <= " 998";
            when 997 => reg0_string <= " 997";
            when 996 => reg0_string <= " 996";
            when 995 => reg0_string <= " 995";
            when 994 => reg0_string <= " 994";
            when 993 => reg0_string <= " 993";
            when 992 => reg0_string <= " 992";
            when 991 => reg0_string <= " 991";
            when 990 => reg0_string <= " 990";
            when 989 => reg0_string <= " 989";
            when 988 => reg0_string <= " 988";
            when 987 => reg0_string <= " 987";
            when 986 => reg0_string <= " 986";
            when 985 => reg0_string <= " 985";
            when 984 => reg0_string <= " 984";
            when 983 => reg0_string <= " 983";
            when 982 => reg0_string <= " 982";
            when 981 => reg0_string <= " 981";
            when 980 => reg0_string <= " 980";
            when 979 => reg0_string <= " 979";
            when 978 => reg0_string <= " 978";
            when 977 => reg0_string <= " 977";
            when 976 => reg0_string <= " 976";
            when 975 => reg0_string <= " 975";
            when 974 => reg0_string <= " 974";
            when 973 => reg0_string <= " 973";
            when 972 => reg0_string <= " 972";
            when 971 => reg0_string <= " 971";
            when 970 => reg0_string <= " 970";
            when 969 => reg0_string <= " 969";
            when 968 => reg0_string <= " 968";
            when 967 => reg0_string <= " 967";
            when 966 => reg0_string <= " 966";
            when 965 => reg0_string <= " 965";
            when 964 => reg0_string <= " 964";
            when 963 => reg0_string <= " 963";
            when 962 => reg0_string <= " 962";
            when 961 => reg0_string <= " 961";
            when 960 => reg0_string <= " 960";
            when 959 => reg0_string <= " 959";
            when 958 => reg0_string <= " 958";
            when 957 => reg0_string <= " 957";
            when 956 => reg0_string <= " 956";
            when 955 => reg0_string <= " 955";
            when 954 => reg0_string <= " 954";
            when 953 => reg0_string <= " 953";
            when 952 => reg0_string <= " 952";
            when 951 => reg0_string <= " 951";
            when 950 => reg0_string <= " 950";
            when 949 => reg0_string <= " 949";
            when 948 => reg0_string <= " 948";
            when 947 => reg0_string <= " 947";
            when 946 => reg0_string <= " 946";
            when 945 => reg0_string <= " 945";
            when 944 => reg0_string <= " 944";
            when 943 => reg0_string <= " 943";
            when 942 => reg0_string <= " 942";
            when 941 => reg0_string <= " 941";
            when 940 => reg0_string <= " 940";
            when 939 => reg0_string <= " 939";
            when 938 => reg0_string <= " 938";
            when 937 => reg0_string <= " 937";
            when 936 => reg0_string <= " 936";
            when 935 => reg0_string <= " 935";
            when 934 => reg0_string <= " 934";
            when 933 => reg0_string <= " 933";
            when 932 => reg0_string <= " 932";
            when 931 => reg0_string <= " 931";
            when 930 => reg0_string <= " 930";
            when 929 => reg0_string <= " 929";
            when 928 => reg0_string <= " 928";
            when 927 => reg0_string <= " 927";
            when 926 => reg0_string <= " 926";
            when 925 => reg0_string <= " 925";
            when 924 => reg0_string <= " 924";
            when 923 => reg0_string <= " 923";
            when 922 => reg0_string <= " 922";
            when 921 => reg0_string <= " 921";
            when 920 => reg0_string <= " 920";
            when 919 => reg0_string <= " 919";
            when 918 => reg0_string <= " 918";
            when 917 => reg0_string <= " 917";
            when 916 => reg0_string <= " 916";
            when 915 => reg0_string <= " 915";
            when 914 => reg0_string <= " 914";
            when 913 => reg0_string <= " 913";
            when 912 => reg0_string <= " 912";
            when 911 => reg0_string <= " 911";
            when 910 => reg0_string <= " 910";
            when 909 => reg0_string <= " 909";
            when 908 => reg0_string <= " 908";
            when 907 => reg0_string <= " 907";
            when 906 => reg0_string <= " 906";
            when 905 => reg0_string <= " 905";
            when 904 => reg0_string <= " 904";
            when 903 => reg0_string <= " 903";
            when 902 => reg0_string <= " 902";
            when 901 => reg0_string <= " 901";
            when 900 => reg0_string <= " 900";
            when 899 => reg0_string <= " 899";
            when 898 => reg0_string <= " 898";
            when 897 => reg0_string <= " 897";
            when 896 => reg0_string <= " 896";
            when 895 => reg0_string <= " 895";
            when 894 => reg0_string <= " 894";
            when 893 => reg0_string <= " 893";
            when 892 => reg0_string <= " 892";
            when 891 => reg0_string <= " 891";
            when 890 => reg0_string <= " 890";
            when 889 => reg0_string <= " 889";
            when 888 => reg0_string <= " 888";
            when 887 => reg0_string <= " 887";
            when 886 => reg0_string <= " 886";
            when 885 => reg0_string <= " 885";
            when 884 => reg0_string <= " 884";
            when 883 => reg0_string <= " 883";
            when 882 => reg0_string <= " 882";
            when 881 => reg0_string <= " 881";
            when 880 => reg0_string <= " 880";
            when 879 => reg0_string <= " 879";
            when 878 => reg0_string <= " 878";
            when 877 => reg0_string <= " 877";
            when 876 => reg0_string <= " 876";
            when 875 => reg0_string <= " 875";
            when 874 => reg0_string <= " 874";
            when 873 => reg0_string <= " 873";
            when 872 => reg0_string <= " 872";
            when 871 => reg0_string <= " 871";
            when 870 => reg0_string <= " 870";
            when 869 => reg0_string <= " 869";
            when 868 => reg0_string <= " 868";
            when 867 => reg0_string <= " 867";
            when 866 => reg0_string <= " 866";
            when 865 => reg0_string <= " 865";
            when 864 => reg0_string <= " 864";
            when 863 => reg0_string <= " 863";
            when 862 => reg0_string <= " 862";
            when 861 => reg0_string <= " 861";
            when 860 => reg0_string <= " 860";
            when 859 => reg0_string <= " 859";
            when 858 => reg0_string <= " 858";
            when 857 => reg0_string <= " 857";
            when 856 => reg0_string <= " 856";
            when 855 => reg0_string <= " 855";
            when 854 => reg0_string <= " 854";
            when 853 => reg0_string <= " 853";
            when 852 => reg0_string <= " 852";
            when 851 => reg0_string <= " 851";
            when 850 => reg0_string <= " 850";
            when 849 => reg0_string <= " 849";
            when 848 => reg0_string <= " 848";
            when 847 => reg0_string <= " 847";
            when 846 => reg0_string <= " 846";
            when 845 => reg0_string <= " 845";
            when 844 => reg0_string <= " 844";
            when 843 => reg0_string <= " 843";
            when 842 => reg0_string <= " 842";
            when 841 => reg0_string <= " 841";
            when 840 => reg0_string <= " 840";
            when 839 => reg0_string <= " 839";
            when 838 => reg0_string <= " 838";
            when 837 => reg0_string <= " 837";
            when 836 => reg0_string <= " 836";
            when 835 => reg0_string <= " 835";
            when 834 => reg0_string <= " 834";
            when 833 => reg0_string <= " 833";
            when 832 => reg0_string <= " 832";
            when 831 => reg0_string <= " 831";
            when 830 => reg0_string <= " 830";
            when 829 => reg0_string <= " 829";
            when 828 => reg0_string <= " 828";
            when 827 => reg0_string <= " 827";
            when 826 => reg0_string <= " 826";
            when 825 => reg0_string <= " 825";
            when 824 => reg0_string <= " 824";
            when 823 => reg0_string <= " 823";
            when 822 => reg0_string <= " 822";
            when 821 => reg0_string <= " 821";
            when 820 => reg0_string <= " 820";
            when 819 => reg0_string <= " 819";
            when 818 => reg0_string <= " 818";
            when 817 => reg0_string <= " 817";
            when 816 => reg0_string <= " 816";
            when 815 => reg0_string <= " 815";
            when 814 => reg0_string <= " 814";
            when 813 => reg0_string <= " 813";
            when 812 => reg0_string <= " 812";
            when 811 => reg0_string <= " 811";
            when 810 => reg0_string <= " 810";
            when 809 => reg0_string <= " 809";
            when 808 => reg0_string <= " 808";
            when 807 => reg0_string <= " 807";
            when 806 => reg0_string <= " 806";
            when 805 => reg0_string <= " 805";
            when 804 => reg0_string <= " 804";
            when 803 => reg0_string <= " 803";
            when 802 => reg0_string <= " 802";
            when 801 => reg0_string <= " 801";
            when 800 => reg0_string <= " 800";
            when 799 => reg0_string <= " 799";
            when 798 => reg0_string <= " 798";
            when 797 => reg0_string <= " 797";
            when 796 => reg0_string <= " 796";
            when 795 => reg0_string <= " 795";
            when 794 => reg0_string <= " 794";
            when 793 => reg0_string <= " 793";
            when 792 => reg0_string <= " 792";
            when 791 => reg0_string <= " 791";
            when 790 => reg0_string <= " 790";
            when 789 => reg0_string <= " 789";
            when 788 => reg0_string <= " 788";
            when 787 => reg0_string <= " 787";
            when 786 => reg0_string <= " 786";
            when 785 => reg0_string <= " 785";
            when 784 => reg0_string <= " 784";
            when 783 => reg0_string <= " 783";
            when 782 => reg0_string <= " 782";
            when 781 => reg0_string <= " 781";
            when 780 => reg0_string <= " 780";
            when 779 => reg0_string <= " 779";
            when 778 => reg0_string <= " 778";
            when 777 => reg0_string <= " 777";
            when 776 => reg0_string <= " 776";
            when 775 => reg0_string <= " 775";
            when 774 => reg0_string <= " 774";
            when 773 => reg0_string <= " 773";
            when 772 => reg0_string <= " 772";
            when 771 => reg0_string <= " 771";
            when 770 => reg0_string <= " 770";
            when 769 => reg0_string <= " 769";
            when 768 => reg0_string <= " 768";
            when 767 => reg0_string <= " 767";
            when 766 => reg0_string <= " 766";
            when 765 => reg0_string <= " 765";
            when 764 => reg0_string <= " 764";
            when 763 => reg0_string <= " 763";
            when 762 => reg0_string <= " 762";
            when 761 => reg0_string <= " 761";
            when 760 => reg0_string <= " 760";
            when 759 => reg0_string <= " 759";
            when 758 => reg0_string <= " 758";
            when 757 => reg0_string <= " 757";
            when 756 => reg0_string <= " 756";
            when 755 => reg0_string <= " 755";
            when 754 => reg0_string <= " 754";
            when 753 => reg0_string <= " 753";
            when 752 => reg0_string <= " 752";
            when 751 => reg0_string <= " 751";
            when 750 => reg0_string <= " 750";
            when 749 => reg0_string <= " 749";
            when 748 => reg0_string <= " 748";
            when 747 => reg0_string <= " 747";
            when 746 => reg0_string <= " 746";
            when 745 => reg0_string <= " 745";
            when 744 => reg0_string <= " 744";
            when 743 => reg0_string <= " 743";
            when 742 => reg0_string <= " 742";
            when 741 => reg0_string <= " 741";
            when 740 => reg0_string <= " 740";
            when 739 => reg0_string <= " 739";
            when 738 => reg0_string <= " 738";
            when 737 => reg0_string <= " 737";
            when 736 => reg0_string <= " 736";
            when 735 => reg0_string <= " 735";
            when 734 => reg0_string <= " 734";
            when 733 => reg0_string <= " 733";
            when 732 => reg0_string <= " 732";
            when 731 => reg0_string <= " 731";
            when 730 => reg0_string <= " 730";
            when 729 => reg0_string <= " 729";
            when 728 => reg0_string <= " 728";
            when 727 => reg0_string <= " 727";
            when 726 => reg0_string <= " 726";
            when 725 => reg0_string <= " 725";
            when 724 => reg0_string <= " 724";
            when 723 => reg0_string <= " 723";
            when 722 => reg0_string <= " 722";
            when 721 => reg0_string <= " 721";
            when 720 => reg0_string <= " 720";
            when 719 => reg0_string <= " 719";
            when 718 => reg0_string <= " 718";
            when 717 => reg0_string <= " 717";
            when 716 => reg0_string <= " 716";
            when 715 => reg0_string <= " 715";
            when 714 => reg0_string <= " 714";
            when 713 => reg0_string <= " 713";
            when 712 => reg0_string <= " 712";
            when 711 => reg0_string <= " 711";
            when 710 => reg0_string <= " 710";
            when 709 => reg0_string <= " 709";
            when 708 => reg0_string <= " 708";
            when 707 => reg0_string <= " 707";
            when 706 => reg0_string <= " 706";
            when 705 => reg0_string <= " 705";
            when 704 => reg0_string <= " 704";
            when 703 => reg0_string <= " 703";
            when 702 => reg0_string <= " 702";
            when 701 => reg0_string <= " 701";
            when 700 => reg0_string <= " 700";
            when 699 => reg0_string <= " 699";
            when 698 => reg0_string <= " 698";
            when 697 => reg0_string <= " 697";
            when 696 => reg0_string <= " 696";
            when 695 => reg0_string <= " 695";
            when 694 => reg0_string <= " 694";
            when 693 => reg0_string <= " 693";
            when 692 => reg0_string <= " 692";
            when 691 => reg0_string <= " 691";
            when 690 => reg0_string <= " 690";
            when 689 => reg0_string <= " 689";
            when 688 => reg0_string <= " 688";
            when 687 => reg0_string <= " 687";
            when 686 => reg0_string <= " 686";
            when 685 => reg0_string <= " 685";
            when 684 => reg0_string <= " 684";
            when 683 => reg0_string <= " 683";
            when 682 => reg0_string <= " 682";
            when 681 => reg0_string <= " 681";
            when 680 => reg0_string <= " 680";
            when 679 => reg0_string <= " 679";
            when 678 => reg0_string <= " 678";
            when 677 => reg0_string <= " 677";
            when 676 => reg0_string <= " 676";
            when 675 => reg0_string <= " 675";
            when 674 => reg0_string <= " 674";
            when 673 => reg0_string <= " 673";
            when 672 => reg0_string <= " 672";
            when 671 => reg0_string <= " 671";
            when 670 => reg0_string <= " 670";
            when 669 => reg0_string <= " 669";
            when 668 => reg0_string <= " 668";
            when 667 => reg0_string <= " 667";
            when 666 => reg0_string <= " 666";
            when 665 => reg0_string <= " 665";
            when 664 => reg0_string <= " 664";
            when 663 => reg0_string <= " 663";
            when 662 => reg0_string <= " 662";
            when 661 => reg0_string <= " 661";
            when 660 => reg0_string <= " 660";
            when 659 => reg0_string <= " 659";
            when 658 => reg0_string <= " 658";
            when 657 => reg0_string <= " 657";
            when 656 => reg0_string <= " 656";
            when 655 => reg0_string <= " 655";
            when 654 => reg0_string <= " 654";
            when 653 => reg0_string <= " 653";
            when 652 => reg0_string <= " 652";
            when 651 => reg0_string <= " 651";
            when 650 => reg0_string <= " 650";
            when 649 => reg0_string <= " 649";
            when 648 => reg0_string <= " 648";
            when 647 => reg0_string <= " 647";
            when 646 => reg0_string <= " 646";
            when 645 => reg0_string <= " 645";
            when 644 => reg0_string <= " 644";
            when 643 => reg0_string <= " 643";
            when 642 => reg0_string <= " 642";
            when 641 => reg0_string <= " 641";
            when 640 => reg0_string <= " 640";
            when 639 => reg0_string <= " 639";
            when 638 => reg0_string <= " 638";
            when 637 => reg0_string <= " 637";
            when 636 => reg0_string <= " 636";
            when 635 => reg0_string <= " 635";
            when 634 => reg0_string <= " 634";
            when 633 => reg0_string <= " 633";
            when 632 => reg0_string <= " 632";
            when 631 => reg0_string <= " 631";
            when 630 => reg0_string <= " 630";
            when 629 => reg0_string <= " 629";
            when 628 => reg0_string <= " 628";
            when 627 => reg0_string <= " 627";
            when 626 => reg0_string <= " 626";
            when 625 => reg0_string <= " 625";
            when 624 => reg0_string <= " 624";
            when 623 => reg0_string <= " 623";
            when 622 => reg0_string <= " 622";
            when 621 => reg0_string <= " 621";
            when 620 => reg0_string <= " 620";
            when 619 => reg0_string <= " 619";
            when 618 => reg0_string <= " 618";
            when 617 => reg0_string <= " 617";
            when 616 => reg0_string <= " 616";
            when 615 => reg0_string <= " 615";
            when 614 => reg0_string <= " 614";
            when 613 => reg0_string <= " 613";
            when 612 => reg0_string <= " 612";
            when 611 => reg0_string <= " 611";
            when 610 => reg0_string <= " 610";
            when 609 => reg0_string <= " 609";
            when 608 => reg0_string <= " 608";
            when 607 => reg0_string <= " 607";
            when 606 => reg0_string <= " 606";
            when 605 => reg0_string <= " 605";
            when 604 => reg0_string <= " 604";
            when 603 => reg0_string <= " 603";
            when 602 => reg0_string <= " 602";
            when 601 => reg0_string <= " 601";
            when 600 => reg0_string <= " 600";
            when 599 => reg0_string <= " 599";
            when 598 => reg0_string <= " 598";
            when 597 => reg0_string <= " 597";
            when 596 => reg0_string <= " 596";
            when 595 => reg0_string <= " 595";
            when 594 => reg0_string <= " 594";
            when 593 => reg0_string <= " 593";
            when 592 => reg0_string <= " 592";
            when 591 => reg0_string <= " 591";
            when 590 => reg0_string <= " 590";
            when 589 => reg0_string <= " 589";
            when 588 => reg0_string <= " 588";
            when 587 => reg0_string <= " 587";
            when 586 => reg0_string <= " 586";
            when 585 => reg0_string <= " 585";
            when 584 => reg0_string <= " 584";
            when 583 => reg0_string <= " 583";
            when 582 => reg0_string <= " 582";
            when 581 => reg0_string <= " 581";
            when 580 => reg0_string <= " 580";
            when 579 => reg0_string <= " 579";
            when 578 => reg0_string <= " 578";
            when 577 => reg0_string <= " 577";
            when 576 => reg0_string <= " 576";
            when 575 => reg0_string <= " 575";
            when 574 => reg0_string <= " 574";
            when 573 => reg0_string <= " 573";
            when 572 => reg0_string <= " 572";
            when 571 => reg0_string <= " 571";
            when 570 => reg0_string <= " 570";
            when 569 => reg0_string <= " 569";
            when 568 => reg0_string <= " 568";
            when 567 => reg0_string <= " 567";
            when 566 => reg0_string <= " 566";
            when 565 => reg0_string <= " 565";
            when 564 => reg0_string <= " 564";
            when 563 => reg0_string <= " 563";
            when 562 => reg0_string <= " 562";
            when 561 => reg0_string <= " 561";
            when 560 => reg0_string <= " 560";
            when 559 => reg0_string <= " 559";
            when 558 => reg0_string <= " 558";
            when 557 => reg0_string <= " 557";
            when 556 => reg0_string <= " 556";
            when 555 => reg0_string <= " 555";
            when 554 => reg0_string <= " 554";
            when 553 => reg0_string <= " 553";
            when 552 => reg0_string <= " 552";
            when 551 => reg0_string <= " 551";
            when 550 => reg0_string <= " 550";
            when 549 => reg0_string <= " 549";
            when 548 => reg0_string <= " 548";
            when 547 => reg0_string <= " 547";
            when 546 => reg0_string <= " 546";
            when 545 => reg0_string <= " 545";
            when 544 => reg0_string <= " 544";
            when 543 => reg0_string <= " 543";
            when 542 => reg0_string <= " 542";
            when 541 => reg0_string <= " 541";
            when 540 => reg0_string <= " 540";
            when 539 => reg0_string <= " 539";
            when 538 => reg0_string <= " 538";
            when 537 => reg0_string <= " 537";
            when 536 => reg0_string <= " 536";
            when 535 => reg0_string <= " 535";
            when 534 => reg0_string <= " 534";
            when 533 => reg0_string <= " 533";
            when 532 => reg0_string <= " 532";
            when 531 => reg0_string <= " 531";
            when 530 => reg0_string <= " 530";
            when 529 => reg0_string <= " 529";
            when 528 => reg0_string <= " 528";
            when 527 => reg0_string <= " 527";
            when 526 => reg0_string <= " 526";
            when 525 => reg0_string <= " 525";
            when 524 => reg0_string <= " 524";
            when 523 => reg0_string <= " 523";
            when 522 => reg0_string <= " 522";
            when 521 => reg0_string <= " 521";
            when 520 => reg0_string <= " 520";
            when 519 => reg0_string <= " 519";
            when 518 => reg0_string <= " 518";
            when 517 => reg0_string <= " 517";
            when 516 => reg0_string <= " 516";
            when 515 => reg0_string <= " 515";
            when 514 => reg0_string <= " 514";
            when 513 => reg0_string <= " 513";
            when 512 => reg0_string <= " 512";
            when 511 => reg0_string <= " 511";
            when 510 => reg0_string <= " 510";
            when 509 => reg0_string <= " 509";
            when 508 => reg0_string <= " 508";
            when 507 => reg0_string <= " 507";
            when 506 => reg0_string <= " 506";
            when 505 => reg0_string <= " 505";
            when 504 => reg0_string <= " 504";
            when 503 => reg0_string <= " 503";
            when 502 => reg0_string <= " 502";
            when 501 => reg0_string <= " 501";
            when 500 => reg0_string <= " 500";
            when 499 => reg0_string <= " 499";
            when 498 => reg0_string <= " 498";
            when 497 => reg0_string <= " 497";
            when 496 => reg0_string <= " 496";
            when 495 => reg0_string <= " 495";
            when 494 => reg0_string <= " 494";
            when 493 => reg0_string <= " 493";
            when 492 => reg0_string <= " 492";
            when 491 => reg0_string <= " 491";
            when 490 => reg0_string <= " 490";
            when 489 => reg0_string <= " 489";
            when 488 => reg0_string <= " 488";
            when 487 => reg0_string <= " 487";
            when 486 => reg0_string <= " 486";
            when 485 => reg0_string <= " 485";
            when 484 => reg0_string <= " 484";
            when 483 => reg0_string <= " 483";
            when 482 => reg0_string <= " 482";
            when 481 => reg0_string <= " 481";
            when 480 => reg0_string <= " 480";
            when 479 => reg0_string <= " 479";
            when 478 => reg0_string <= " 478";
            when 477 => reg0_string <= " 477";
            when 476 => reg0_string <= " 476";
            when 475 => reg0_string <= " 475";
            when 474 => reg0_string <= " 474";
            when 473 => reg0_string <= " 473";
            when 472 => reg0_string <= " 472";
            when 471 => reg0_string <= " 471";
            when 470 => reg0_string <= " 470";
            when 469 => reg0_string <= " 469";
            when 468 => reg0_string <= " 468";
            when 467 => reg0_string <= " 467";
            when 466 => reg0_string <= " 466";
            when 465 => reg0_string <= " 465";
            when 464 => reg0_string <= " 464";
            when 463 => reg0_string <= " 463";
            when 462 => reg0_string <= " 462";
            when 461 => reg0_string <= " 461";
            when 460 => reg0_string <= " 460";
            when 459 => reg0_string <= " 459";
            when 458 => reg0_string <= " 458";
            when 457 => reg0_string <= " 457";
            when 456 => reg0_string <= " 456";
            when 455 => reg0_string <= " 455";
            when 454 => reg0_string <= " 454";
            when 453 => reg0_string <= " 453";
            when 452 => reg0_string <= " 452";
            when 451 => reg0_string <= " 451";
            when 450 => reg0_string <= " 450";
            when 449 => reg0_string <= " 449";
            when 448 => reg0_string <= " 448";
            when 447 => reg0_string <= " 447";
            when 446 => reg0_string <= " 446";
            when 445 => reg0_string <= " 445";
            when 444 => reg0_string <= " 444";
            when 443 => reg0_string <= " 443";
            when 442 => reg0_string <= " 442";
            when 441 => reg0_string <= " 441";
            when 440 => reg0_string <= " 440";
            when 439 => reg0_string <= " 439";
            when 438 => reg0_string <= " 438";
            when 437 => reg0_string <= " 437";
            when 436 => reg0_string <= " 436";
            when 435 => reg0_string <= " 435";
            when 434 => reg0_string <= " 434";
            when 433 => reg0_string <= " 433";
            when 432 => reg0_string <= " 432";
            when 431 => reg0_string <= " 431";
            when 430 => reg0_string <= " 430";
            when 429 => reg0_string <= " 429";
            when 428 => reg0_string <= " 428";
            when 427 => reg0_string <= " 427";
            when 426 => reg0_string <= " 426";
            when 425 => reg0_string <= " 425";
            when 424 => reg0_string <= " 424";
            when 423 => reg0_string <= " 423";
            when 422 => reg0_string <= " 422";
            when 421 => reg0_string <= " 421";
            when 420 => reg0_string <= " 420";
            when 419 => reg0_string <= " 419";
            when 418 => reg0_string <= " 418";
            when 417 => reg0_string <= " 417";
            when 416 => reg0_string <= " 416";
            when 415 => reg0_string <= " 415";
            when 414 => reg0_string <= " 414";
            when 413 => reg0_string <= " 413";
            when 412 => reg0_string <= " 412";
            when 411 => reg0_string <= " 411";
            when 410 => reg0_string <= " 410";
            when 409 => reg0_string <= " 409";
            when 408 => reg0_string <= " 408";
            when 407 => reg0_string <= " 407";
            when 406 => reg0_string <= " 406";
            when 405 => reg0_string <= " 405";
            when 404 => reg0_string <= " 404";
            when 403 => reg0_string <= " 403";
            when 402 => reg0_string <= " 402";
            when 401 => reg0_string <= " 401";
            when 400 => reg0_string <= " 400";
            when 399 => reg0_string <= " 399";
            when 398 => reg0_string <= " 398";
            when 397 => reg0_string <= " 397";
            when 396 => reg0_string <= " 396";
            when 395 => reg0_string <= " 395";
            when 394 => reg0_string <= " 394";
            when 393 => reg0_string <= " 393";
            when 392 => reg0_string <= " 392";
            when 391 => reg0_string <= " 391";
            when 390 => reg0_string <= " 390";
            when 389 => reg0_string <= " 389";
            when 388 => reg0_string <= " 388";
            when 387 => reg0_string <= " 387";
            when 386 => reg0_string <= " 386";
            when 385 => reg0_string <= " 385";
            when 384 => reg0_string <= " 384";
            when 383 => reg0_string <= " 383";
            when 382 => reg0_string <= " 382";
            when 381 => reg0_string <= " 381";
            when 380 => reg0_string <= " 380";
            when 379 => reg0_string <= " 379";
            when 378 => reg0_string <= " 378";
            when 377 => reg0_string <= " 377";
            when 376 => reg0_string <= " 376";
            when 375 => reg0_string <= " 375";
            when 374 => reg0_string <= " 374";
            when 373 => reg0_string <= " 373";
            when 372 => reg0_string <= " 372";
            when 371 => reg0_string <= " 371";
            when 370 => reg0_string <= " 370";
            when 369 => reg0_string <= " 369";
            when 368 => reg0_string <= " 368";
            when 367 => reg0_string <= " 367";
            when 366 => reg0_string <= " 366";
            when 365 => reg0_string <= " 365";
            when 364 => reg0_string <= " 364";
            when 363 => reg0_string <= " 363";
            when 362 => reg0_string <= " 362";
            when 361 => reg0_string <= " 361";
            when 360 => reg0_string <= " 360";
            when 359 => reg0_string <= " 359";
            when 358 => reg0_string <= " 358";
            when 357 => reg0_string <= " 357";
            when 356 => reg0_string <= " 356";
            when 355 => reg0_string <= " 355";
            when 354 => reg0_string <= " 354";
            when 353 => reg0_string <= " 353";
            when 352 => reg0_string <= " 352";
            when 351 => reg0_string <= " 351";
            when 350 => reg0_string <= " 350";
            when 349 => reg0_string <= " 349";
            when 348 => reg0_string <= " 348";
            when 347 => reg0_string <= " 347";
            when 346 => reg0_string <= " 346";
            when 345 => reg0_string <= " 345";
            when 344 => reg0_string <= " 344";
            when 343 => reg0_string <= " 343";
            when 342 => reg0_string <= " 342";
            when 341 => reg0_string <= " 341";
            when 340 => reg0_string <= " 340";
            when 339 => reg0_string <= " 339";
            when 338 => reg0_string <= " 338";
            when 337 => reg0_string <= " 337";
            when 336 => reg0_string <= " 336";
            when 335 => reg0_string <= " 335";
            when 334 => reg0_string <= " 334";
            when 333 => reg0_string <= " 333";
            when 332 => reg0_string <= " 332";
            when 331 => reg0_string <= " 331";
            when 330 => reg0_string <= " 330";
            when 329 => reg0_string <= " 329";
            when 328 => reg0_string <= " 328";
            when 327 => reg0_string <= " 327";
            when 326 => reg0_string <= " 326";
            when 325 => reg0_string <= " 325";
            when 324 => reg0_string <= " 324";
            when 323 => reg0_string <= " 323";
            when 322 => reg0_string <= " 322";
            when 321 => reg0_string <= " 321";
            when 320 => reg0_string <= " 320";
            when 319 => reg0_string <= " 319";
            when 318 => reg0_string <= " 318";
            when 317 => reg0_string <= " 317";
            when 316 => reg0_string <= " 316";
            when 315 => reg0_string <= " 315";
            when 314 => reg0_string <= " 314";
            when 313 => reg0_string <= " 313";
            when 312 => reg0_string <= " 312";
            when 311 => reg0_string <= " 311";
            when 310 => reg0_string <= " 310";
            when 309 => reg0_string <= " 309";
            when 308 => reg0_string <= " 308";
            when 307 => reg0_string <= " 307";
            when 306 => reg0_string <= " 306";
            when 305 => reg0_string <= " 305";
            when 304 => reg0_string <= " 304";
            when 303 => reg0_string <= " 303";
            when 302 => reg0_string <= " 302";
            when 301 => reg0_string <= " 301";
            when 300 => reg0_string <= " 300";
            when 299 => reg0_string <= " 299";
            when 298 => reg0_string <= " 298";
            when 297 => reg0_string <= " 297";
            when 296 => reg0_string <= " 296";
            when 295 => reg0_string <= " 295";
            when 294 => reg0_string <= " 294";
            when 293 => reg0_string <= " 293";
            when 292 => reg0_string <= " 292";
            when 291 => reg0_string <= " 291";
            when 290 => reg0_string <= " 290";
            when 289 => reg0_string <= " 289";
            when 288 => reg0_string <= " 288";
            when 287 => reg0_string <= " 287";
            when 286 => reg0_string <= " 286";
            when 285 => reg0_string <= " 285";
            when 284 => reg0_string <= " 284";
            when 283 => reg0_string <= " 283";
            when 282 => reg0_string <= " 282";
            when 281 => reg0_string <= " 281";
            when 280 => reg0_string <= " 280";
            when 279 => reg0_string <= " 279";
            when 278 => reg0_string <= " 278";
            when 277 => reg0_string <= " 277";
            when 276 => reg0_string <= " 276";
            when 275 => reg0_string <= " 275";
            when 274 => reg0_string <= " 274";
            when 273 => reg0_string <= " 273";
            when 272 => reg0_string <= " 272";
            when 271 => reg0_string <= " 271";
            when 270 => reg0_string <= " 270";
            when 269 => reg0_string <= " 269";
            when 268 => reg0_string <= " 268";
            when 267 => reg0_string <= " 267";
            when 266 => reg0_string <= " 266";
            when 265 => reg0_string <= " 265";
            when 264 => reg0_string <= " 264";
            when 263 => reg0_string <= " 263";
            when 262 => reg0_string <= " 262";
            when 261 => reg0_string <= " 261";
            when 260 => reg0_string <= " 260";
            when 259 => reg0_string <= " 259";
            when 258 => reg0_string <= " 258";
            when 257 => reg0_string <= " 257";
            when 256 => reg0_string <= " 256";
            when 255 => reg0_string <= " 255";
            when 254 => reg0_string <= " 254";
            when 253 => reg0_string <= " 253";
            when 252 => reg0_string <= " 252";
            when 251 => reg0_string <= " 251";
            when 250 => reg0_string <= " 250";
            when 249 => reg0_string <= " 249";
            when 248 => reg0_string <= " 248";
            when 247 => reg0_string <= " 247";
            when 246 => reg0_string <= " 246";
            when 245 => reg0_string <= " 245";
            when 244 => reg0_string <= " 244";
            when 243 => reg0_string <= " 243";
            when 242 => reg0_string <= " 242";
            when 241 => reg0_string <= " 241";
            when 240 => reg0_string <= " 240";
            when 239 => reg0_string <= " 239";
            when 238 => reg0_string <= " 238";
            when 237 => reg0_string <= " 237";
            when 236 => reg0_string <= " 236";
            when 235 => reg0_string <= " 235";
            when 234 => reg0_string <= " 234";
            when 233 => reg0_string <= " 233";
            when 232 => reg0_string <= " 232";
            when 231 => reg0_string <= " 231";
            when 230 => reg0_string <= " 230";
            when 229 => reg0_string <= " 229";
            when 228 => reg0_string <= " 228";
            when 227 => reg0_string <= " 227";
            when 226 => reg0_string <= " 226";
            when 225 => reg0_string <= " 225";
            when 224 => reg0_string <= " 224";
            when 223 => reg0_string <= " 223";
            when 222 => reg0_string <= " 222";
            when 221 => reg0_string <= " 221";
            when 220 => reg0_string <= " 220";
            when 219 => reg0_string <= " 219";
            when 218 => reg0_string <= " 218";
            when 217 => reg0_string <= " 217";
            when 216 => reg0_string <= " 216";
            when 215 => reg0_string <= " 215";
            when 214 => reg0_string <= " 214";
            when 213 => reg0_string <= " 213";
            when 212 => reg0_string <= " 212";
            when 211 => reg0_string <= " 211";
            when 210 => reg0_string <= " 210";
            when 209 => reg0_string <= " 209";
            when 208 => reg0_string <= " 208";
            when 207 => reg0_string <= " 207";
            when 206 => reg0_string <= " 206";
            when 205 => reg0_string <= " 205";
            when 204 => reg0_string <= " 204";
            when 203 => reg0_string <= " 203";
            when 202 => reg0_string <= " 202";
            when 201 => reg0_string <= " 201";
            when 200 => reg0_string <= " 200";
            when 199 => reg0_string <= " 199";
            when 198 => reg0_string <= " 198";
            when 197 => reg0_string <= " 197";
            when 196 => reg0_string <= " 196";
            when 195 => reg0_string <= " 195";
            when 194 => reg0_string <= " 194";
            when 193 => reg0_string <= " 193";
            when 192 => reg0_string <= " 192";
            when 191 => reg0_string <= " 191";
            when 190 => reg0_string <= " 190";
            when 189 => reg0_string <= " 189";
            when 188 => reg0_string <= " 188";
            when 187 => reg0_string <= " 187";
            when 186 => reg0_string <= " 186";
            when 185 => reg0_string <= " 185";
            when 184 => reg0_string <= " 184";
            when 183 => reg0_string <= " 183";
            when 182 => reg0_string <= " 182";
            when 181 => reg0_string <= " 181";
            when 180 => reg0_string <= " 180";
            when 179 => reg0_string <= " 179";
            when 178 => reg0_string <= " 178";
            when 177 => reg0_string <= " 177";
            when 176 => reg0_string <= " 176";
            when 175 => reg0_string <= " 175";
            when 174 => reg0_string <= " 174";
            when 173 => reg0_string <= " 173";
            when 172 => reg0_string <= " 172";
            when 171 => reg0_string <= " 171";
            when 170 => reg0_string <= " 170";
            when 169 => reg0_string <= " 169";
            when 168 => reg0_string <= " 168";
            when 167 => reg0_string <= " 167";
            when 166 => reg0_string <= " 166";
            when 165 => reg0_string <= " 165";
            when 164 => reg0_string <= " 164";
            when 163 => reg0_string <= " 163";
            when 162 => reg0_string <= " 162";
            when 161 => reg0_string <= " 161";
            when 160 => reg0_string <= " 160";
            when 159 => reg0_string <= " 159";
            when 158 => reg0_string <= " 158";
            when 157 => reg0_string <= " 157";
            when 156 => reg0_string <= " 156";
            when 155 => reg0_string <= " 155";
            when 154 => reg0_string <= " 154";
            when 153 => reg0_string <= " 153";
            when 152 => reg0_string <= " 152";
            when 151 => reg0_string <= " 151";
            when 150 => reg0_string <= " 150";
            when 149 => reg0_string <= " 149";
            when 148 => reg0_string <= " 148";
            when 147 => reg0_string <= " 147";
            when 146 => reg0_string <= " 146";
            when 145 => reg0_string <= " 145";
            when 144 => reg0_string <= " 144";
            when 143 => reg0_string <= " 143";
            when 142 => reg0_string <= " 142";
            when 141 => reg0_string <= " 141";
            when 140 => reg0_string <= " 140";
            when 139 => reg0_string <= " 139";
            when 138 => reg0_string <= " 138";
            when 137 => reg0_string <= " 137";
            when 136 => reg0_string <= " 136";
            when 135 => reg0_string <= " 135";
            when 134 => reg0_string <= " 134";
            when 133 => reg0_string <= " 133";
            when 132 => reg0_string <= " 132";
            when 131 => reg0_string <= " 131";
            when 130 => reg0_string <= " 130";
            when 129 => reg0_string <= " 129";
            when 128 => reg0_string <= " 128";
            when 127 => reg0_string <= " 127";
            when 126 => reg0_string <= " 126";
            when 125 => reg0_string <= " 125";
            when 124 => reg0_string <= " 124";
            when 123 => reg0_string <= " 123";
            when 122 => reg0_string <= " 122";
            when 121 => reg0_string <= " 121";
            when 120 => reg0_string <= " 120";
            when 119 => reg0_string <= " 119";
            when 118 => reg0_string <= " 118";
            when 117 => reg0_string <= " 117";
            when 116 => reg0_string <= " 116";
            when 115 => reg0_string <= " 115";
            when 114 => reg0_string <= " 114";
            when 113 => reg0_string <= " 113";
            when 112 => reg0_string <= " 112";
            when 111 => reg0_string <= " 111";
            when 110 => reg0_string <= " 110";
            when 109 => reg0_string <= " 109";
            when 108 => reg0_string <= " 108";
            when 107 => reg0_string <= " 107";                                                                                        
            when 106 => reg0_string <= " 106";                                                                                        
            when 105 => reg0_string <= " 105";                                                                                        
            when 104 => reg0_string <= " 104";                                                                                        
            when 103 => reg0_string <= " 103";                                                                                        
            when 102 => reg0_string <= " 102";                                                                                        
            when 101 => reg0_string <= " 101";                                                                                        
            when 100 => reg0_string <= " 100";                                                                                        
            when 99 => reg0_string <= "  99";                                                                                         
            when 98 => reg0_string <= "  98";                                                                                         
            when 97 => reg0_string <= "  97";                                                                                         
            when 96 => reg0_string <= "  96";                                                                                         
            when 95 => reg0_string <= "  95";                                                                                         
            when 94 => reg0_string <= "  94";                                                                                         
            when 93 => reg0_string <= "  93";                                                                                         
            when 92 => reg0_string <= "  92";                                                                                         
            when 91 => reg0_string <= "  91";                                                                                         
            when 90 => reg0_string <= "  90";                                                                                         
            when 89 => reg0_string <= "  89";                                                                                         
            when 88 => reg0_string <= "  88";                                                                                         
            when 87 => reg0_string <= "  87";                                                                                         
            when 86 => reg0_string <= "  86";                                                                                         
            when 85 => reg0_string <= "  85";                                                                                         
            when 84 => reg0_string <= "  84";                                                                                         
            when 83 => reg0_string <= "  83";                                                                                         
            when 82 => reg0_string <= "  82";                                                                                         
            when 81 => reg0_string <= "  81";                                                                                         
            when 80 => reg0_string <= "  80";                                                                                         
            when 79 => reg0_string <= "  79";                                                                                         
            when 78 => reg0_string <= "  78";                                                                                         
            when 77 => reg0_string <= "  77";
            when 76 => reg0_string <= "  76";                                                                                         
            when 75 => reg0_string <= "  75";                                                                                         
            when 74 => reg0_string <= "  74";                                                                                         
            when 73 => reg0_string <= "  73";                                                                                         
            when 72 => reg0_string <= "  72";                                                                                         
            when 71 => reg0_string <= "  71";                                                                                         
            when 70 => reg0_string <= "  70";                                                                                         
            when 69 => reg0_string <= "  69";                                                                                         
            when 68 => reg0_string <= "  68";                                                                                         
            when 67 => reg0_string <= "  67";                                                                                         
            when 66 => reg0_string <= "  66";                                                                                         
            when 65 => reg0_string <= "  65";                                                                                         
            when 64 => reg0_string <= "  64";                                                                                         
            when 63 => reg0_string <= "  63";                                                                                         
            when 62 => reg0_string <= "  62";                                                                                         
            when 61 => reg0_string <= "  61";                                                                                         
            when 60 => reg0_string <= "  60";                                                                                         
            when 59 => reg0_string <= "  59";                                                                                         
            when 58 => reg0_string <= "  58";                                                                                         
            when 57 => reg0_string <= "  57";                                                                                         
            when 56 => reg0_string <= "  56";                                                                                         
            when 55 => reg0_string <= "  55";                                                                                         
            when 54 => reg0_string <= "  54";                                                                                         
            when 53 => reg0_string <= "  53";                                                                                         
            when 52 => reg0_string <= "  52";                                                                                         
            when 51 => reg0_string <= "  51";                                                                                         
            when 50 => reg0_string <= "  50";                                                                                         
            when 49 => reg0_string <= "  49";                                                                                         
            when 48 => reg0_string <= "  48";                                                                                         
            when 47 => reg0_string <= "  47";
            when 46 => reg0_string <= "  46";                                                                                         
            when 45 => reg0_string <= "  45";                                                                                         
            when 44 => reg0_string <= "  44";                                                                                         
            when 43 => reg0_string <= "  43";                                                                                         
            when 42 => reg0_string <= "  42";                                                                                         
            when 41 => reg0_string <= "  41";                                                                                         
            when 40 => reg0_string <= "  40";                                                                                         
            when 39 => reg0_string <= "  39";                                                                                         
            when 38 => reg0_string <= "  38";                                                                                         
            when 37 => reg0_string <= "  37";                                                                                         
            when 36 => reg0_string <= "  36";                                                                                         
            when 35 => reg0_string <= "  35";                                                                                         
            when 34 => reg0_string <= "  34";                                                                                         
            when 33 => reg0_string <= "  33";                                                                                         
            when 32 => reg0_string <= "  32";                                                                                         
            when 31 => reg0_string <= "  31";                                                                                         
            when 30 => reg0_string <= "  30";                                                                                         
            when 29 => reg0_string <= "  29";                                                                                         
            when 28 => reg0_string <= "  28";                                                                                         
            when 27 => reg0_string <= "  27";                                                                                         
            when 26 => reg0_string <= "  26";                                                                                         
            when 25 => reg0_string <= "  25";                                                                                         
            when 24 => reg0_string <= "  24";                                                                                         
            when 23 => reg0_string <= "  23";
            when 22 => reg0_string <= "  22";                                                                                         
            when 21 => reg0_string <= "  21";                                                                                         
            when 20 => reg0_string <= "  20";                                                                                         
            when 19 => reg0_string <= "  19";                                                                                         
            when 18 => reg0_string <= "  18";                                                                                         
            when 17 => reg0_string <= "  17";                                                                                         
            when 16 => reg0_string <= "  16";                                                                                         
            when 15 => reg0_string <= "  15";                                                                                         
            when 14 => reg0_string <= "  14";                                                                                         
            when 13 => reg0_string <= "  13";                                                                                         
            when 12 => reg0_string <= "  12";                                                                                         
            when 11 => reg0_string <= "  11";                                                                                         
            when 10 => reg0_string <= "  10";                                                                                         
            when 9  => reg0_string <= "   9";                                                                                          
            when 8  => reg0_string <= "   8";                                                                                          
            when 7  => reg0_string <= "   7";                                                                                          
            when 6  => reg0_string <= "   6";                                                                                          
            when 5  => reg0_string <= "   5";                                                                                          
            when 4  => reg0_string <= "   4";                                                                                          
            when 3  => reg0_string <= "   3";                                                                                          
            when 2  => reg0_string <= "   2";                                                                                          
            when 1  => reg0_string <= "   1";                                                                                          
            when 0  => reg0_string <= "   0";
            when -1 => reg0_string <= "  -1";
            when -2 => reg0_string <= "  -2";
            when -3 => reg0_string <= "  -3";
            when -4 => reg0_string <= "  -4";
            when -5 => reg0_string <= "  -5";
            when -6 => reg0_string <= "  -6";
            when -7 => reg0_string <= "  -7";
            when -8 => reg0_string <= "  -8";
            when -9 => reg0_string <= "  -9";
            when -10 => reg0_string <= " -10";
            when -11 => reg0_string <= " -11";
            when -12 => reg0_string <= " -12";
            when -13 => reg0_string <= " -13";
            when -14 => reg0_string <= " -14";
            when -15 => reg0_string <= " -15";
            when -16 => reg0_string <= " -16";
            when -17 => reg0_string <= " -17";
            when -18 => reg0_string <= " -18";
            when -19 => reg0_string <= " -19";
            when -20 => reg0_string <= " -20";
            when -21 => reg0_string <= " -21";
            when -22 => reg0_string <= " -22";
            when -23 => reg0_string <= " -23";
            when -24 => reg0_string <= " -24";
            when -25 => reg0_string <= " -25";
            when -26 => reg0_string <= " -26";
            when -27 => reg0_string <= " -27";
            when -28 => reg0_string <= " -28";
            when -29 => reg0_string <= " -29";
            when -30 => reg0_string <= " -30";
            when -31 => reg0_string <= " -31";
            when -32 => reg0_string <= " -32";
            when -33 => reg0_string <= " -33";
            when -34 => reg0_string <= " -34";
            when -35 => reg0_string <= " -35";
            when -36 => reg0_string <= " -36";
            when -37 => reg0_string <= " -37";
            when -38 => reg0_string <= " -38";
            when -39 => reg0_string <= " -39";
            when -40 => reg0_string <= " -40";
            when -41 => reg0_string <= " -41";
            when -42 => reg0_string <= " -42";
            when -43 => reg0_string <= " -43";
            when -44 => reg0_string <= " -44";
            when -45 => reg0_string <= " -45";
            when -46 => reg0_string <= " -46";
            when -47 => reg0_string <= " -47";
            when -48 => reg0_string <= " -48";
            when -49 => reg0_string <= " -49";
            when -50 => reg0_string <= " -50";
            when -51 => reg0_string <= " -51";
            when -52 => reg0_string <= " -52";
            when -53 => reg0_string <= " -53";
            when -54 => reg0_string <= " -54";
            when -55 => reg0_string <= " -55";
            when -56 => reg0_string <= " -56";
            when -57 => reg0_string <= " -57";
            when -58 => reg0_string <= " -58";
            when -59 => reg0_string <= " -59";
            when -60 => reg0_string <= " -60";
            when -61 => reg0_string <= " -61";
            when -62 => reg0_string <= " -62";
            when -63 => reg0_string <= " -63";
            when -64 => reg0_string <= " -64";
            when -65 => reg0_string <= " -65";
            when -66 => reg0_string <= " -66";
            when -67 => reg0_string <= " -67";
            when -68 => reg0_string <= " -68";
            when -69 => reg0_string <= " -69";
            when -70 => reg0_string <= " -70";
            when -71 => reg0_string <= " -71";
            when -72 => reg0_string <= " -72";
            when -73 => reg0_string <= " -73";
            when -74 => reg0_string <= " -74";
            when -75 => reg0_string <= " -75";
            when -76 => reg0_string <= " -76";
            when -77 => reg0_string <= " -77";
            when -78 => reg0_string <= " -78";
            when -79 => reg0_string <= " -79";
            when -80 => reg0_string <= " -80";
            when -81 => reg0_string <= " -81";
            when -82 => reg0_string <= " -82";
            when -83 => reg0_string <= " -83";
            when -84 => reg0_string <= " -84";
            when -85 => reg0_string <= " -85";
            when -86 => reg0_string <= " -86";
            when -87 => reg0_string <= " -87";
            when -88 => reg0_string <= " -88";
            when -89 => reg0_string <= " -89";
            when -90 => reg0_string <= " -90";
            when -91 => reg0_string <= " -91";
            when -92 => reg0_string <= " -92";
            when -93 => reg0_string <= " -93";
            when -94 => reg0_string <= " -94";
            when -95 => reg0_string <= " -95";
            when -96 => reg0_string <= " -96";
            when -97 => reg0_string <= " -97";
            when -98 => reg0_string <= " -98";
            when -99 => reg0_string <= " -99";
            when -100 => reg0_string <= "-100";
            when -101 => reg0_string <= "-101";
            when -102 => reg0_string <= "-102";
            when -103 => reg0_string <= "-103";
            when -104 => reg0_string <= "-104";
            when -105 => reg0_string <= "-105";
            when -106 => reg0_string <= "-106";
            when -107 => reg0_string <= "-107";
            when -108 => reg0_string <= "-108";
            when -109 => reg0_string <= "-109";
            when -110 => reg0_string <= "-110";
            when -111 => reg0_string <= "-111";
            when -112 => reg0_string <= "-112";
            when -113 => reg0_string <= "-113";
            when -114 => reg0_string <= "-114";
            when -115 => reg0_string <= "-115";
            when -116 => reg0_string <= "-116";
            when -117 => reg0_string <= "-117";
            when -118 => reg0_string <= "-118";
            when -119 => reg0_string <= "-119";
            when -120 => reg0_string <= "-120";
            when -121 => reg0_string <= "-121";
            when -122 => reg0_string <= "-122";
            when -123 => reg0_string <= "-123";
            when -124 => reg0_string <= "-124";
            when -125 => reg0_string <= "-125";
            when -126 => reg0_string <= "-126";
            when -127 => reg0_string <= "-127";
            when -128 => reg0_string <= "-128";
            when -129 => reg0_string <= "-129";
            when -130 => reg0_string <= "-130";
            when -131 => reg0_string <= "-131";
            when -132 => reg0_string <= "-132";
            when -133 => reg0_string <= "-133";
            when -134 => reg0_string <= "-134";
            when -135 => reg0_string <= "-135";
            when -136 => reg0_string <= "-136";
            when -137 => reg0_string <= "-137";
            when -138 => reg0_string <= "-138";
            when -139 => reg0_string <= "-139";
            when -140 => reg0_string <= "-140";
            when -141 => reg0_string <= "-141";
            when -142 => reg0_string <= "-142";
            when -143 => reg0_string <= "-143";
            when -144 => reg0_string <= "-144";
            when -145 => reg0_string <= "-145";
            when -146 => reg0_string <= "-146";
            when -147 => reg0_string <= "-147";
            when -148 => reg0_string <= "-148";
            when -149 => reg0_string <= "-149";
            when -150 => reg0_string <= "-150";
            when -151 => reg0_string <= "-151";
            when -152 => reg0_string <= "-152";
            when -153 => reg0_string <= "-153";
            when -154 => reg0_string <= "-154";
            when -155 => reg0_string <= "-155";
            when -156 => reg0_string <= "-156";
            when -157 => reg0_string <= "-157";
            when -158 => reg0_string <= "-158";
            when -159 => reg0_string <= "-159";
            when -160 => reg0_string <= "-160";
            when -161 => reg0_string <= "-161";
            when -162 => reg0_string <= "-162";
            when -163 => reg0_string <= "-163";
            when -164 => reg0_string <= "-164";
            when -165 => reg0_string <= "-165";
            when -166 => reg0_string <= "-166";
            when -167 => reg0_string <= "-167";
            when -168 => reg0_string <= "-168";
            when -169 => reg0_string <= "-169";
            when -170 => reg0_string <= "-170";
            when -171 => reg0_string <= "-171";
            when -172 => reg0_string <= "-172";
            when -173 => reg0_string <= "-173";
            when -174 => reg0_string <= "-174";
            when -175 => reg0_string <= "-175";
            when -176 => reg0_string <= "-176";
            when -177 => reg0_string <= "-177";
            when -178 => reg0_string <= "-178";
            when -179 => reg0_string <= "-179";
            when -180 => reg0_string <= "-180";
            when -181 => reg0_string <= "-181";
            when -182 => reg0_string <= "-182";
            when -183 => reg0_string <= "-183";
            when -184 => reg0_string <= "-184";
            when -185 => reg0_string <= "-185";
            when -186 => reg0_string <= "-186";
            when -187 => reg0_string <= "-187";
            when -188 => reg0_string <= "-188";
            when -189 => reg0_string <= "-189";
            when -190 => reg0_string <= "-190";
            when -191 => reg0_string <= "-191";
            when -192 => reg0_string <= "-192";
            when -193 => reg0_string <= "-193";
            when -194 => reg0_string <= "-194";
            when -195 => reg0_string <= "-195";
            when -196 => reg0_string <= "-196";
            when -197 => reg0_string <= "-197";
            when -198 => reg0_string <= "-198";
            when -199 => reg0_string <= "-199";
            when -200 => reg0_string <= "-200";
            when -201 => reg0_string <= "-201";
            when -202 => reg0_string <= "-202";
            when -203 => reg0_string <= "-203";
            when -204 => reg0_string <= "-204";
            when -205 => reg0_string <= "-205";
            when -206 => reg0_string <= "-206";
            when -207 => reg0_string <= "-207";
            when -208 => reg0_string <= "-208";
            when -209 => reg0_string <= "-209";
            when -210 => reg0_string <= "-210";
            when -211 => reg0_string <= "-211";
            when -212 => reg0_string <= "-212";
            when -213 => reg0_string <= "-213";
            when -214 => reg0_string <= "-214";
            when -215 => reg0_string <= "-215";
            when -216 => reg0_string <= "-216";
            when -217 => reg0_string <= "-217";
            when -218 => reg0_string <= "-218";
            when -219 => reg0_string <= "-219";
            when -220 => reg0_string <= "-220";
            when -221 => reg0_string <= "-221";
            when -222 => reg0_string <= "-222";
            when -223 => reg0_string <= "-223";
            when -224 => reg0_string <= "-224";
            when -225 => reg0_string <= "-225";
            when -226 => reg0_string <= "-226";
            when -227 => reg0_string <= "-227";
            when -228 => reg0_string <= "-228";
            when -229 => reg0_string <= "-229";
            when -230 => reg0_string <= "-230";
            when -231 => reg0_string <= "-231";
            when -232 => reg0_string <= "-232";
            when -233 => reg0_string <= "-233";
            when -234 => reg0_string <= "-234";
            when -235 => reg0_string <= "-235";
            when -236 => reg0_string <= "-236";
            when -237 => reg0_string <= "-237";
            when -238 => reg0_string <= "-238";
            when -239 => reg0_string <= "-239";
            when -240 => reg0_string <= "-240";
            when -241 => reg0_string <= "-241";
            when -242 => reg0_string <= "-242";
            when -243 => reg0_string <= "-243";
            when -244 => reg0_string <= "-244";
            when -245 => reg0_string <= "-245";
            when -246 => reg0_string <= "-246";
            when -247 => reg0_string <= "-247";
            when -248 => reg0_string <= "-248";
            when -249 => reg0_string <= "-249";
            when -250 => reg0_string <= "-250";
            when -251 => reg0_string <= "-251";
            when -252 => reg0_string <= "-252";
            when -253 => reg0_string <= "-253";
            when -254 => reg0_string <= "-254";
            when -255 => reg0_string <= "-255";
            when -256 => reg0_string <= "-256";
            when -257 => reg0_string <= "-257";
            when -258 => reg0_string <= "-258";
            when -259 => reg0_string <= "-259";
            when -260 => reg0_string <= "-260";
            when -261 => reg0_string <= "-261";
            when -262 => reg0_string <= "-262";
            when -263 => reg0_string <= "-263";
            when -264 => reg0_string <= "-264";
            when -265 => reg0_string <= "-265";
            when -266 => reg0_string <= "-266";
            when -267 => reg0_string <= "-267";
            when -268 => reg0_string <= "-268";
            when -269 => reg0_string <= "-269";
            when -270 => reg0_string <= "-270";
            when -271 => reg0_string <= "-271";
            when -272 => reg0_string <= "-272";
            when -273 => reg0_string <= "-273";
            when -274 => reg0_string <= "-274";
            when -275 => reg0_string <= "-275";
            when -276 => reg0_string <= "-276";
            when -277 => reg0_string <= "-277";
            when -278 => reg0_string <= "-278";
            when -279 => reg0_string <= "-279";
            when -280 => reg0_string <= "-280";
            when -281 => reg0_string <= "-281";
            when -282 => reg0_string <= "-282";
            when -283 => reg0_string <= "-283";
            when -284 => reg0_string <= "-284";
            when -285 => reg0_string <= "-285";
            when -286 => reg0_string <= "-286";
            when -287 => reg0_string <= "-287";
            when -288 => reg0_string <= "-288";
            when -289 => reg0_string <= "-289";
            when -290 => reg0_string <= "-290";
            when -291 => reg0_string <= "-291";
            when -292 => reg0_string <= "-292";
            when -293 => reg0_string <= "-293";
            when -294 => reg0_string <= "-294";
            when -295 => reg0_string <= "-295";
            when -296 => reg0_string <= "-296";
            when -297 => reg0_string <= "-297";
            when -298 => reg0_string <= "-298";
            when -299 => reg0_string <= "-299";
            when -300 => reg0_string <= "-300";
            when -301 => reg0_string <= "-301";
            when -302 => reg0_string <= "-302";
            when -303 => reg0_string <= "-303";
            when -304 => reg0_string <= "-304";
            when -305 => reg0_string <= "-305";
            when -306 => reg0_string <= "-306";
            when -307 => reg0_string <= "-307";
            when -308 => reg0_string <= "-308";
            when -309 => reg0_string <= "-309";
            when -310 => reg0_string <= "-310";
            when -311 => reg0_string <= "-311";
            when -312 => reg0_string <= "-312";
            when -313 => reg0_string <= "-313";
            when -314 => reg0_string <= "-314";
            when -315 => reg0_string <= "-315";
            when -316 => reg0_string <= "-316";
            when -317 => reg0_string <= "-317";
            when -318 => reg0_string <= "-318";
            when -319 => reg0_string <= "-319";
            when -320 => reg0_string <= "-320";
            when -321 => reg0_string <= "-321";
            when -322 => reg0_string <= "-322";
            when -323 => reg0_string <= "-323";
            when -324 => reg0_string <= "-324";
            when -325 => reg0_string <= "-325";
            when -326 => reg0_string <= "-326";
            when -327 => reg0_string <= "-327";
            when -328 => reg0_string <= "-328";
            when -329 => reg0_string <= "-329";
            when -330 => reg0_string <= "-330";
            when -331 => reg0_string <= "-331";
            when -332 => reg0_string <= "-332";
            when -333 => reg0_string <= "-333";
            when -334 => reg0_string <= "-334";
            when -335 => reg0_string <= "-335";
            when -336 => reg0_string <= "-336";
            when -337 => reg0_string <= "-337";
            when -338 => reg0_string <= "-338";
            when -339 => reg0_string <= "-339";
            when -340 => reg0_string <= "-340";
            when -341 => reg0_string <= "-341";
            when -342 => reg0_string <= "-342";
            when -343 => reg0_string <= "-343";
            when -344 => reg0_string <= "-344";
            when -345 => reg0_string <= "-345";
            when -346 => reg0_string <= "-346";
            when -347 => reg0_string <= "-347";
            when -348 => reg0_string <= "-348";
            when -349 => reg0_string <= "-349";
            when -350 => reg0_string <= "-350";
            when -351 => reg0_string <= "-351";
            when -352 => reg0_string <= "-352";
            when -353 => reg0_string <= "-353";
            when -354 => reg0_string <= "-354";
            when -355 => reg0_string <= "-355";
            when -356 => reg0_string <= "-356";
            when -357 => reg0_string <= "-357";
            when -358 => reg0_string <= "-358";
            when -359 => reg0_string <= "-359";
            when -360 => reg0_string <= "-360";
            when -361 => reg0_string <= "-361";
            when -362 => reg0_string <= "-362";
            when -363 => reg0_string <= "-363";
            when -364 => reg0_string <= "-364";
            when -365 => reg0_string <= "-365";
            when -366 => reg0_string <= "-366";
            when -367 => reg0_string <= "-367";
            when -368 => reg0_string <= "-368";
            when -369 => reg0_string <= "-369";
            when -370 => reg0_string <= "-370";
            when -371 => reg0_string <= "-371";
            when -372 => reg0_string <= "-372";
            when -373 => reg0_string <= "-373";
            when -374 => reg0_string <= "-374";
            when -375 => reg0_string <= "-375";
            when -376 => reg0_string <= "-376";
            when -377 => reg0_string <= "-377";
            when -378 => reg0_string <= "-378";
            when -379 => reg0_string <= "-379";
            when -380 => reg0_string <= "-380";
            when -381 => reg0_string <= "-381";
            when -382 => reg0_string <= "-382";
            when -383 => reg0_string <= "-383";
            when -384 => reg0_string <= "-384";
            when -385 => reg0_string <= "-385";
            when -386 => reg0_string <= "-386";
            when -387 => reg0_string <= "-387";
            when -388 => reg0_string <= "-388";
            when -389 => reg0_string <= "-389";
            when -390 => reg0_string <= "-390";
            when -391 => reg0_string <= "-391";
            when -392 => reg0_string <= "-392";
            when -393 => reg0_string <= "-393";
            when -394 => reg0_string <= "-394";
            when -395 => reg0_string <= "-395";
            when -396 => reg0_string <= "-396";
            when -397 => reg0_string <= "-397";
            when -398 => reg0_string <= "-398";
            when -399 => reg0_string <= "-399";
            when -400 => reg0_string <= "-400";
            when -401 => reg0_string <= "-401";
            when -402 => reg0_string <= "-402";
            when -403 => reg0_string <= "-403";
            when -404 => reg0_string <= "-404";
            when -405 => reg0_string <= "-405";
            when -406 => reg0_string <= "-406";
            when -407 => reg0_string <= "-407";
            when -408 => reg0_string <= "-408";
            when -409 => reg0_string <= "-409";
            when -410 => reg0_string <= "-410";
            when -411 => reg0_string <= "-411";
            when -412 => reg0_string <= "-412";
            when -413 => reg0_string <= "-413";
            when -414 => reg0_string <= "-414";
            when -415 => reg0_string <= "-415";
            when -416 => reg0_string <= "-416";
            when -417 => reg0_string <= "-417";
            when -418 => reg0_string <= "-418";
            when -419 => reg0_string <= "-419";
            when -420 => reg0_string <= "-420";
            when -421 => reg0_string <= "-421";
            when -422 => reg0_string <= "-422";
            when -423 => reg0_string <= "-423";
            when -424 => reg0_string <= "-424";
            when -425 => reg0_string <= "-425";
            when -426 => reg0_string <= "-426";
            when -427 => reg0_string <= "-427";
            when -428 => reg0_string <= "-428";
            when -429 => reg0_string <= "-429";
            when -430 => reg0_string <= "-430";
            when -431 => reg0_string <= "-431";
            when -432 => reg0_string <= "-432";
            when -433 => reg0_string <= "-433";
            when -434 => reg0_string <= "-434";
            when -435 => reg0_string <= "-435";
            when -436 => reg0_string <= "-436";
            when -437 => reg0_string <= "-437";
            when -438 => reg0_string <= "-438";
            when -439 => reg0_string <= "-439";
            when -440 => reg0_string <= "-440";
            when -441 => reg0_string <= "-441";
            when -442 => reg0_string <= "-442";
            when -443 => reg0_string <= "-443";
            when -444 => reg0_string <= "-444";
            when -445 => reg0_string <= "-445";
            when -446 => reg0_string <= "-446";
            when -447 => reg0_string <= "-447";
            when -448 => reg0_string <= "-448";
            when -449 => reg0_string <= "-449";
            when -450 => reg0_string <= "-450";
            when -451 => reg0_string <= "-451";
            when -452 => reg0_string <= "-452";
            when -453 => reg0_string <= "-453";
            when -454 => reg0_string <= "-454";
            when -455 => reg0_string <= "-455";
            when -456 => reg0_string <= "-456";
            when -457 => reg0_string <= "-457";
            when -458 => reg0_string <= "-458";
            when -459 => reg0_string <= "-459";
            when -460 => reg0_string <= "-460";
            when -461 => reg0_string <= "-461";
            when -462 => reg0_string <= "-462";
            when -463 => reg0_string <= "-463";
            when -464 => reg0_string <= "-464";
            when -465 => reg0_string <= "-465";
            when -466 => reg0_string <= "-466";
            when -467 => reg0_string <= "-467";
            when -468 => reg0_string <= "-468";
            when -469 => reg0_string <= "-469";
            when -470 => reg0_string <= "-470";
            when -471 => reg0_string <= "-471";
            when -472 => reg0_string <= "-472";
            when -473 => reg0_string <= "-473";
            when -474 => reg0_string <= "-474";
            when -475 => reg0_string <= "-475";
            when -476 => reg0_string <= "-476";
            when -477 => reg0_string <= "-477";
            when -478 => reg0_string <= "-478";
            when -479 => reg0_string <= "-479";
            when -480 => reg0_string <= "-480";
            when -481 => reg0_string <= "-481";
            when -482 => reg0_string <= "-482";
            when -483 => reg0_string <= "-483";
            when -484 => reg0_string <= "-484";
            when -485 => reg0_string <= "-485";
            when -486 => reg0_string <= "-486";
            when -487 => reg0_string <= "-487";
            when -488 => reg0_string <= "-488";
            when -489 => reg0_string <= "-489";
            when -490 => reg0_string <= "-490";
            when -491 => reg0_string <= "-491";
            when -492 => reg0_string <= "-492";
            when -493 => reg0_string <= "-493";
            when -494 => reg0_string <= "-494";
            when -495 => reg0_string <= "-495";
            when -496 => reg0_string <= "-496";
            when -497 => reg0_string <= "-497";
            when -498 => reg0_string <= "-498";
            when -499 => reg0_string <= "-499";
            when -500 => reg0_string <= "-500";
            when -501 => reg0_string <= "-501";
            when -502 => reg0_string <= "-502";
            when -503 => reg0_string <= "-503";
            when -504 => reg0_string <= "-504";
            when -505 => reg0_string <= "-505";
            when -506 => reg0_string <= "-506";
            when -507 => reg0_string <= "-507";
            when -508 => reg0_string <= "-508";
            when -509 => reg0_string <= "-509";
            when -510 => reg0_string <= "-510";
            when -511 => reg0_string <= "-511";
            when -512 => reg0_string <= "-512";
            when -513 => reg0_string <= "-513";
            when -514 => reg0_string <= "-514";
            when -515 => reg0_string <= "-515";
            when -516 => reg0_string <= "-516";
            when -517 => reg0_string <= "-517";
            when -518 => reg0_string <= "-518";
            when -519 => reg0_string <= "-519";
            when -520 => reg0_string <= "-520";
            when -521 => reg0_string <= "-521";
            when -522 => reg0_string <= "-522";
            when -523 => reg0_string <= "-523";
            when -524 => reg0_string <= "-524";
            when -525 => reg0_string <= "-525";
            when -526 => reg0_string <= "-526";
            when -527 => reg0_string <= "-527";
            when -528 => reg0_string <= "-528";
            when -529 => reg0_string <= "-529";
            when -530 => reg0_string <= "-530";
            when -531 => reg0_string <= "-531";
            when -532 => reg0_string <= "-532";
            when -533 => reg0_string <= "-533";
            when -534 => reg0_string <= "-534";
            when -535 => reg0_string <= "-535";
            when -536 => reg0_string <= "-536";
            when -537 => reg0_string <= "-537";
            when -538 => reg0_string <= "-538";
            when -539 => reg0_string <= "-539";
            when -540 => reg0_string <= "-540";
            when -541 => reg0_string <= "-541";
            when -542 => reg0_string <= "-542";
            when -543 => reg0_string <= "-543";
            when -544 => reg0_string <= "-544";
            when -545 => reg0_string <= "-545";
            when -546 => reg0_string <= "-546";
            when -547 => reg0_string <= "-547";
            when -548 => reg0_string <= "-548";
            when -549 => reg0_string <= "-549";
            when -550 => reg0_string <= "-550";
            when -551 => reg0_string <= "-551";
            when -552 => reg0_string <= "-552";
            when -553 => reg0_string <= "-553";
            when -554 => reg0_string <= "-554";
            when -555 => reg0_string <= "-555";
            when -556 => reg0_string <= "-556";
            when -557 => reg0_string <= "-557";
            when -558 => reg0_string <= "-558";
            when -559 => reg0_string <= "-559";
            when -560 => reg0_string <= "-560";
            when -561 => reg0_string <= "-561";
            when -562 => reg0_string <= "-562";
            when -563 => reg0_string <= "-563";
            when -564 => reg0_string <= "-564";
            when -565 => reg0_string <= "-565";
            when -566 => reg0_string <= "-566";
            when -567 => reg0_string <= "-567";
            when -568 => reg0_string <= "-568";
            when -569 => reg0_string <= "-569";
            when -570 => reg0_string <= "-570";
            when -571 => reg0_string <= "-571";
            when -572 => reg0_string <= "-572";
            when -573 => reg0_string <= "-573";
            when -574 => reg0_string <= "-574";
            when -575 => reg0_string <= "-575";
            when -576 => reg0_string <= "-576";
            when -577 => reg0_string <= "-577";
            when -578 => reg0_string <= "-578";
            when -579 => reg0_string <= "-579";
            when -580 => reg0_string <= "-580";
            when -581 => reg0_string <= "-581";
            when -582 => reg0_string <= "-582";
            when -583 => reg0_string <= "-583";
            when -584 => reg0_string <= "-584";
            when -585 => reg0_string <= "-585";
            when -586 => reg0_string <= "-586";
            when -587 => reg0_string <= "-587";
            when -588 => reg0_string <= "-588";
            when -589 => reg0_string <= "-589";
            when -590 => reg0_string <= "-590";
            when -591 => reg0_string <= "-591";
            when -592 => reg0_string <= "-592";
            when -593 => reg0_string <= "-593";
            when -594 => reg0_string <= "-594";
            when -595 => reg0_string <= "-595";
            when -596 => reg0_string <= "-596";
            when -597 => reg0_string <= "-597";
            when -598 => reg0_string <= "-598";
            when -599 => reg0_string <= "-599";
            when -600 => reg0_string <= "-600";
            when -601 => reg0_string <= "-601";
            when -602 => reg0_string <= "-602";
            when -603 => reg0_string <= "-603";
            when -604 => reg0_string <= "-604";
            when -605 => reg0_string <= "-605";
            when -606 => reg0_string <= "-606";
            when -607 => reg0_string <= "-607";
            when -608 => reg0_string <= "-608";
            when -609 => reg0_string <= "-609";
            when -610 => reg0_string <= "-610";
            when -611 => reg0_string <= "-611";
            when -612 => reg0_string <= "-612";
            when -613 => reg0_string <= "-613";
            when -614 => reg0_string <= "-614";
            when -615 => reg0_string <= "-615";
            when -616 => reg0_string <= "-616";
            when -617 => reg0_string <= "-617";
            when -618 => reg0_string <= "-618";
            when -619 => reg0_string <= "-619";
            when -620 => reg0_string <= "-620";
            when -621 => reg0_string <= "-621";
            when -622 => reg0_string <= "-622";
            when -623 => reg0_string <= "-623";
            when -624 => reg0_string <= "-624";
            when -625 => reg0_string <= "-625";
            when -626 => reg0_string <= "-626";
            when -627 => reg0_string <= "-627";
            when -628 => reg0_string <= "-628";
            when -629 => reg0_string <= "-629";
            when -630 => reg0_string <= "-630";
            when -631 => reg0_string <= "-631";
            when -632 => reg0_string <= "-632";
            when -633 => reg0_string <= "-633";
            when -634 => reg0_string <= "-634";
            when -635 => reg0_string <= "-635";
            when -636 => reg0_string <= "-636";
            when -637 => reg0_string <= "-637";
            when -638 => reg0_string <= "-638";
            when -639 => reg0_string <= "-639";
            when -640 => reg0_string <= "-640";
            when -641 => reg0_string <= "-641";
            when -642 => reg0_string <= "-642";
            when -643 => reg0_string <= "-643";
            when -644 => reg0_string <= "-644";
            when -645 => reg0_string <= "-645";
            when -646 => reg0_string <= "-646";
            when -647 => reg0_string <= "-647";
            when -648 => reg0_string <= "-648";
            when -649 => reg0_string <= "-649";
            when -650 => reg0_string <= "-650";
            when -651 => reg0_string <= "-651";
            when -652 => reg0_string <= "-652";
            when -653 => reg0_string <= "-653";
            when -654 => reg0_string <= "-654";
            when -655 => reg0_string <= "-655";
            when -656 => reg0_string <= "-656";
            when -657 => reg0_string <= "-657";
            when -658 => reg0_string <= "-658";
            when -659 => reg0_string <= "-659";
            when -660 => reg0_string <= "-660";
            when -661 => reg0_string <= "-661";
            when -662 => reg0_string <= "-662";
            when -663 => reg0_string <= "-663";
            when -664 => reg0_string <= "-664";
            when -665 => reg0_string <= "-665";
            when -666 => reg0_string <= "-666";
            when -667 => reg0_string <= "-667";
            when -668 => reg0_string <= "-668";
            when -669 => reg0_string <= "-669";
            when -670 => reg0_string <= "-670";
            when -671 => reg0_string <= "-671";
            when -672 => reg0_string <= "-672";
            when -673 => reg0_string <= "-673";
            when -674 => reg0_string <= "-674";
            when -675 => reg0_string <= "-675";
            when -676 => reg0_string <= "-676";
            when -677 => reg0_string <= "-677";
            when -678 => reg0_string <= "-678";
            when -679 => reg0_string <= "-679";
            when -680 => reg0_string <= "-680";
            when -681 => reg0_string <= "-681";
            when -682 => reg0_string <= "-682";
            when -683 => reg0_string <= "-683";
            when -684 => reg0_string <= "-684";
            when -685 => reg0_string <= "-685";
            when -686 => reg0_string <= "-686";
            when -687 => reg0_string <= "-687";
            when -688 => reg0_string <= "-688";
            when -689 => reg0_string <= "-689";
            when -690 => reg0_string <= "-690";
            when -691 => reg0_string <= "-691";
            when -692 => reg0_string <= "-692";
            when -693 => reg0_string <= "-693";
            when -694 => reg0_string <= "-694";
            when -695 => reg0_string <= "-695";
            when -696 => reg0_string <= "-696";
            when -697 => reg0_string <= "-697";
            when -698 => reg0_string <= "-698";
            when -699 => reg0_string <= "-699";
            when -700 => reg0_string <= "-700";
            when -701 => reg0_string <= "-701";
            when -702 => reg0_string <= "-702";
            when -703 => reg0_string <= "-703";
            when -704 => reg0_string <= "-704";
            when -705 => reg0_string <= "-705";
            when -706 => reg0_string <= "-706";
            when -707 => reg0_string <= "-707";
            when -708 => reg0_string <= "-708";
            when -709 => reg0_string <= "-709";
            when -710 => reg0_string <= "-710";
            when -711 => reg0_string <= "-711";
            when -712 => reg0_string <= "-712";
            when -713 => reg0_string <= "-713";
            when -714 => reg0_string <= "-714";
            when -715 => reg0_string <= "-715";
            when -716 => reg0_string <= "-716";
            when -717 => reg0_string <= "-717";
            when -718 => reg0_string <= "-718";
            when -719 => reg0_string <= "-719";
            when -720 => reg0_string <= "-720";
            when -721 => reg0_string <= "-721";
            when -722 => reg0_string <= "-722";
            when -723 => reg0_string <= "-723";
            when -724 => reg0_string <= "-724";
            when -725 => reg0_string <= "-725";
            when -726 => reg0_string <= "-726";
            when -727 => reg0_string <= "-727";
            when -728 => reg0_string <= "-728";
            when -729 => reg0_string <= "-729";
            when -730 => reg0_string <= "-730";
            when -731 => reg0_string <= "-731";
            when -732 => reg0_string <= "-732";
            when -733 => reg0_string <= "-733";
            when -734 => reg0_string <= "-734";
            when -735 => reg0_string <= "-735";
            when -736 => reg0_string <= "-736";
            when -737 => reg0_string <= "-737";
            when -738 => reg0_string <= "-738";
            when -739 => reg0_string <= "-739";
            when -740 => reg0_string <= "-740";
            when -741 => reg0_string <= "-741";
            when -742 => reg0_string <= "-742";
            when -743 => reg0_string <= "-743";
            when -744 => reg0_string <= "-744";
            when -745 => reg0_string <= "-745";
            when -746 => reg0_string <= "-746";
            when -747 => reg0_string <= "-747";
            when -748 => reg0_string <= "-748";
            when -749 => reg0_string <= "-749";
            when -750 => reg0_string <= "-750";
            when -751 => reg0_string <= "-751";
            when -752 => reg0_string <= "-752";
            when -753 => reg0_string <= "-753";
            when -754 => reg0_string <= "-754";
            when -755 => reg0_string <= "-755";
            when -756 => reg0_string <= "-756";
            when -757 => reg0_string <= "-757";
            when -758 => reg0_string <= "-758";
            when -759 => reg0_string <= "-759";
            when -760 => reg0_string <= "-760";
            when -761 => reg0_string <= "-761";
            when -762 => reg0_string <= "-762";
            when -763 => reg0_string <= "-763";
            when -764 => reg0_string <= "-764";
            when -765 => reg0_string <= "-765";
            when -766 => reg0_string <= "-766";
            when -767 => reg0_string <= "-767";
            when -768 => reg0_string <= "-768";
            when -769 => reg0_string <= "-769";
            when -770 => reg0_string <= "-770";
            when -771 => reg0_string <= "-771";
            when -772 => reg0_string <= "-772";
            when -773 => reg0_string <= "-773";
            when -774 => reg0_string <= "-774";
            when -775 => reg0_string <= "-775";
            when -776 => reg0_string <= "-776";
            when -777 => reg0_string <= "-777";
            when -778 => reg0_string <= "-778";
            when -779 => reg0_string <= "-779";
            when -780 => reg0_string <= "-780";
            when -781 => reg0_string <= "-781";
            when -782 => reg0_string <= "-782";
            when -783 => reg0_string <= "-783";
            when -784 => reg0_string <= "-784";
            when -785 => reg0_string <= "-785";
            when -786 => reg0_string <= "-786";
            when -787 => reg0_string <= "-787";
            when -788 => reg0_string <= "-788";
            when -789 => reg0_string <= "-789";
            when -790 => reg0_string <= "-790";
            when -791 => reg0_string <= "-791";
            when -792 => reg0_string <= "-792";
            when -793 => reg0_string <= "-793";
            when -794 => reg0_string <= "-794";
            when -795 => reg0_string <= "-795";
            when -796 => reg0_string <= "-796";
            when -797 => reg0_string <= "-797";
            when -798 => reg0_string <= "-798";
            when -799 => reg0_string <= "-799";
            when -800 => reg0_string <= "-800";
            when -801 => reg0_string <= "-801";
            when -802 => reg0_string <= "-802";
            when -803 => reg0_string <= "-803";
            when -804 => reg0_string <= "-804";
            when -805 => reg0_string <= "-805";
            when -806 => reg0_string <= "-806";
            when -807 => reg0_string <= "-807";
            when -808 => reg0_string <= "-808";
            when -809 => reg0_string <= "-809";
            when -810 => reg0_string <= "-810";
            when -811 => reg0_string <= "-811";
            when -812 => reg0_string <= "-812";
            when -813 => reg0_string <= "-813";
            when -814 => reg0_string <= "-814";
            when -815 => reg0_string <= "-815";
            when -816 => reg0_string <= "-816";
            when -817 => reg0_string <= "-817";
            when -818 => reg0_string <= "-818";
            when -819 => reg0_string <= "-819";
            when -820 => reg0_string <= "-820";
            when -821 => reg0_string <= "-821";
            when -822 => reg0_string <= "-822";
            when -823 => reg0_string <= "-823";
            when -824 => reg0_string <= "-824";
            when -825 => reg0_string <= "-825";
            when -826 => reg0_string <= "-826";
            when -827 => reg0_string <= "-827";
            when -828 => reg0_string <= "-828";
            when -829 => reg0_string <= "-829";
            when -830 => reg0_string <= "-830";
            when -831 => reg0_string <= "-831";
            when -832 => reg0_string <= "-832";
            when -833 => reg0_string <= "-833";
            when -834 => reg0_string <= "-834";
            when -835 => reg0_string <= "-835";
            when -836 => reg0_string <= "-836";
            when -837 => reg0_string <= "-837";
            when -838 => reg0_string <= "-838";
            when -839 => reg0_string <= "-839";
            when -840 => reg0_string <= "-840";
            when -841 => reg0_string <= "-841";
            when -842 => reg0_string <= "-842";
            when -843 => reg0_string <= "-843";
            when -844 => reg0_string <= "-844";
            when -845 => reg0_string <= "-845";
            when -846 => reg0_string <= "-846";
            when -847 => reg0_string <= "-847";
            when -848 => reg0_string <= "-848";
            when -849 => reg0_string <= "-849";
            when -850 => reg0_string <= "-850";
            when -851 => reg0_string <= "-851";
            when -852 => reg0_string <= "-852";
            when -853 => reg0_string <= "-853";
            when -854 => reg0_string <= "-854";
            when -855 => reg0_string <= "-855";
            when -856 => reg0_string <= "-856";
            when -857 => reg0_string <= "-857";
            when -858 => reg0_string <= "-858";
            when -859 => reg0_string <= "-859";
            when -860 => reg0_string <= "-860";
            when -861 => reg0_string <= "-861";
            when -862 => reg0_string <= "-862";
            when -863 => reg0_string <= "-863";
            when -864 => reg0_string <= "-864";
            when -865 => reg0_string <= "-865";
            when -866 => reg0_string <= "-866";
            when -867 => reg0_string <= "-867";
            when -868 => reg0_string <= "-868";
            when -869 => reg0_string <= "-869";
            when -870 => reg0_string <= "-870";
            when -871 => reg0_string <= "-871";
            when -872 => reg0_string <= "-872";
            when -873 => reg0_string <= "-873";
            when -874 => reg0_string <= "-874";
            when -875 => reg0_string <= "-875";
            when -876 => reg0_string <= "-876";
            when -877 => reg0_string <= "-877";
            when -878 => reg0_string <= "-878";
            when -879 => reg0_string <= "-879";
            when -880 => reg0_string <= "-880";
            when -881 => reg0_string <= "-881";
            when -882 => reg0_string <= "-882";
            when -883 => reg0_string <= "-883";
            when -884 => reg0_string <= "-884";
            when -885 => reg0_string <= "-885";
            when -886 => reg0_string <= "-886";
            when -887 => reg0_string <= "-887";
            when -888 => reg0_string <= "-888";
            when -889 => reg0_string <= "-889";
            when -890 => reg0_string <= "-890";
            when -891 => reg0_string <= "-891";
            when -892 => reg0_string <= "-892";
            when -893 => reg0_string <= "-893";
            when -894 => reg0_string <= "-894";
            when -895 => reg0_string <= "-895";
            when -896 => reg0_string <= "-896";
            when -897 => reg0_string <= "-897";
            when -898 => reg0_string <= "-898";
            when -899 => reg0_string <= "-899";
            when -900 => reg0_string <= "-900";
            when -901 => reg0_string <= "-901";
            when -902 => reg0_string <= "-902";
            when -903 => reg0_string <= "-903";
            when -904 => reg0_string <= "-904";
            when -905 => reg0_string <= "-905";
            when -906 => reg0_string <= "-906";
            when -907 => reg0_string <= "-907";
            when -908 => reg0_string <= "-908";
            when -909 => reg0_string <= "-909";
            when -910 => reg0_string <= "-910";
            when -911 => reg0_string <= "-911";
            when -912 => reg0_string <= "-912";
            when -913 => reg0_string <= "-913";
            when -914 => reg0_string <= "-914";
            when -915 => reg0_string <= "-915";
            when -916 => reg0_string <= "-916";
            when -917 => reg0_string <= "-917";
            when -918 => reg0_string <= "-918";
            when -919 => reg0_string <= "-919";
            when -920 => reg0_string <= "-920";
            when -921 => reg0_string <= "-921";
            when -922 => reg0_string <= "-922";
            when -923 => reg0_string <= "-923";
            when -924 => reg0_string <= "-924";
            when -925 => reg0_string <= "-925";
            when -926 => reg0_string <= "-926";
            when -927 => reg0_string <= "-927";
            when -928 => reg0_string <= "-928";
            when -929 => reg0_string <= "-929";
            when -930 => reg0_string <= "-930";
            when -931 => reg0_string <= "-931";
            when -932 => reg0_string <= "-932";
            when -933 => reg0_string <= "-933";
            when -934 => reg0_string <= "-934";
            when -935 => reg0_string <= "-935";
            when -936 => reg0_string <= "-936";
            when -937 => reg0_string <= "-937";
            when -938 => reg0_string <= "-938";
            when -939 => reg0_string <= "-939";
            when -940 => reg0_string <= "-940";
            when -941 => reg0_string <= "-941";
            when -942 => reg0_string <= "-942";
            when -943 => reg0_string <= "-943";
            when -944 => reg0_string <= "-944";
            when -945 => reg0_string <= "-945";
            when -946 => reg0_string <= "-946";
            when -947 => reg0_string <= "-947";
            when -948 => reg0_string <= "-948";
            when -949 => reg0_string <= "-949";
            when -950 => reg0_string <= "-950";
            when -951 => reg0_string <= "-951";
            when -952 => reg0_string <= "-952";
            when -953 => reg0_string <= "-953";
            when -954 => reg0_string <= "-954";
            when -955 => reg0_string <= "-955";
            when -956 => reg0_string <= "-956";
            when -957 => reg0_string <= "-957";
            when -958 => reg0_string <= "-958";
            when -959 => reg0_string <= "-959";
            when -960 => reg0_string <= "-960";
            when -961 => reg0_string <= "-961";
            when -962 => reg0_string <= "-962";
            when -963 => reg0_string <= "-963";
            when -964 => reg0_string <= "-964";
            when -965 => reg0_string <= "-965";
            when -966 => reg0_string <= "-966";
            when -967 => reg0_string <= "-967";
            when -968 => reg0_string <= "-968";
            when -969 => reg0_string <= "-969";
            when -970 => reg0_string <= "-970";
            when -971 => reg0_string <= "-971";
            when -972 => reg0_string <= "-972";
            when -973 => reg0_string <= "-973";
            when -974 => reg0_string <= "-974";
            when -975 => reg0_string <= "-975";
            when -976 => reg0_string <= "-976";
            when -977 => reg0_string <= "-977";
            when -978 => reg0_string <= "-978";
            when -979 => reg0_string <= "-979";
            when -980 => reg0_string <= "-980";
            when -981 => reg0_string <= "-981";
            when -982 => reg0_string <= "-982";
            when -983 => reg0_string <= "-983";
            when -984 => reg0_string <= "-984";
            when -985 => reg0_string <= "-985";
            when -986 => reg0_string <= "-986";
            when -987 => reg0_string <= "-987";
            when -988 => reg0_string <= "-988";
            when -989 => reg0_string <= "-989";
            when -990 => reg0_string <= "-990";
            when -991 => reg0_string <= "-991";
            when -992 => reg0_string <= "-992";
            when -993 => reg0_string <= "-993";
            when -994 => reg0_string <= "-994";
            when -995 => reg0_string <= "-995";
            when -996 => reg0_string <= "-996";
            when -997 => reg0_string <= "-997";
            when -998 => reg0_string <= "-998";
            when -999 => reg0_string <= "-999";
            when others => reg0_string <= "    ";
        end case;
    end process;

end Behavioral;
